-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba4",
     9 => x"c0080b0b",
    10 => x"0ba4c408",
    11 => x"0b0b0ba4",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a4c80c0b",
    16 => x"0b0ba4c4",
    17 => x"0c0b0b0b",
    18 => x"a4c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba2b4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a4c070aa",
    57 => x"a0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8fd60402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752e80c7",
    65 => x"38875472",
    66 => x"9c2a7384",
    67 => x"2b545271",
    68 => x"802e8338",
    69 => x"81558972",
    70 => x"259938b7",
    71 => x"1252749b",
    72 => x"38ff1454",
    73 => x"738025df",
    74 => x"38800ba4",
    75 => x"c00c0294",
    76 => x"050d04b0",
    77 => x"12527480",
    78 => x"2ee73871",
    79 => x"5182da2d",
    80 => x"ff145473",
    81 => x"8025c038",
    82 => x"82a904b0",
    83 => x"5182da2d",
    84 => x"800ba4c0",
    85 => x"0c029405",
    86 => x"0d0402f8",
    87 => x"050d7352",
    88 => x"c0087088",
    89 => x"2a708106",
    90 => x"51515170",
    91 => x"802ef138",
    92 => x"71c00c71",
    93 => x"a4c00c02",
    94 => x"88050d04",
    95 => x"02f8050d",
    96 => x"7352c408",
    97 => x"70882a70",
    98 => x"81065151",
    99 => x"5170802e",
   100 => x"f13871c4",
   101 => x"0c71a4c0",
   102 => x"0c028805",
   103 => x"0d0402e8",
   104 => x"050d8078",
   105 => x"57557570",
   106 => x"84055708",
   107 => x"53805472",
   108 => x"982a7388",
   109 => x"2b545271",
   110 => x"802ea238",
   111 => x"c0087088",
   112 => x"2a708106",
   113 => x"51515170",
   114 => x"802ef138",
   115 => x"71c00c81",
   116 => x"15811555",
   117 => x"55837425",
   118 => x"d63871ca",
   119 => x"3874a4c0",
   120 => x"0c029805",
   121 => x"0d0402f4",
   122 => x"050dd452",
   123 => x"81ff720c",
   124 => x"71085381",
   125 => x"ff720c72",
   126 => x"882b83fe",
   127 => x"80067208",
   128 => x"7081ff06",
   129 => x"51525381",
   130 => x"ff720c72",
   131 => x"7107882b",
   132 => x"72087081",
   133 => x"ff065152",
   134 => x"5381ff72",
   135 => x"0c727107",
   136 => x"882b7208",
   137 => x"7081ff06",
   138 => x"7207a4c0",
   139 => x"0c525302",
   140 => x"8c050d04",
   141 => x"02f4050d",
   142 => x"74767181",
   143 => x"ff06d40c",
   144 => x"5353a5a4",
   145 => x"08853871",
   146 => x"892b5271",
   147 => x"982ad40c",
   148 => x"71902a70",
   149 => x"81ff06d4",
   150 => x"0c517188",
   151 => x"2a7081ff",
   152 => x"06d40c51",
   153 => x"7181ff06",
   154 => x"d40c7290",
   155 => x"2a7081ff",
   156 => x"06d40c51",
   157 => x"d4087081",
   158 => x"ff065151",
   159 => x"82b8bf52",
   160 => x"7081ff2e",
   161 => x"09810694",
   162 => x"3881ff0b",
   163 => x"d40cd408",
   164 => x"7081ff06",
   165 => x"ff145451",
   166 => x"5171e538",
   167 => x"70a4c00c",
   168 => x"028c050d",
   169 => x"0402fc05",
   170 => x"0d81c751",
   171 => x"81ff0bd4",
   172 => x"0cff1151",
   173 => x"708025f4",
   174 => x"38028405",
   175 => x"0d0402f0",
   176 => x"050d85a5",
   177 => x"2d819c9f",
   178 => x"53805287",
   179 => x"fc80f751",
   180 => x"84b42da4",
   181 => x"c00854a4",
   182 => x"c008812e",
   183 => x"9038ff13",
   184 => x"5372e638",
   185 => x"72a4c00c",
   186 => x"0290050d",
   187 => x"0481ff0b",
   188 => x"d40c820a",
   189 => x"52849c80",
   190 => x"e95184b4",
   191 => x"2da4c008",
   192 => x"802e8e38",
   193 => x"85a52dff",
   194 => x"135372ff",
   195 => x"bc3885e4",
   196 => x"0481ff0b",
   197 => x"d40c73a4",
   198 => x"c00c0290",
   199 => x"050d0402",
   200 => x"f4050d81",
   201 => x"ff0bd40c",
   202 => x"a2c45183",
   203 => x"9e2d9353",
   204 => x"805287fc",
   205 => x"80c15184",
   206 => x"b42da4c0",
   207 => x"08802e93",
   208 => x"3885a52d",
   209 => x"ff135372",
   210 => x"e73872a4",
   211 => x"c00c028c",
   212 => x"050d0481",
   213 => x"ff0bd40c",
   214 => x"810ba4c0",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050d85a5",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"5184b42d",
   221 => x"a4c00881",
   222 => x"2e8f3886",
   223 => x"9f2d8054",
   224 => x"73a4c00c",
   225 => x"0290050d",
   226 => x"0483e62d",
   227 => x"a4c00883",
   228 => x"ffff0653",
   229 => x"7283aa2e",
   230 => x"098106df",
   231 => x"3881ff0b",
   232 => x"d40cb153",
   233 => x"85be2da4",
   234 => x"c0089538",
   235 => x"72822ece",
   236 => x"38ff1353",
   237 => x"72ee3872",
   238 => x"a4c00c02",
   239 => x"90050d04",
   240 => x"805287fc",
   241 => x"80fa5184",
   242 => x"b42da4c0",
   243 => x"08de3881",
   244 => x"ff0bd40c",
   245 => x"d4085381",
   246 => x"ff0bd40c",
   247 => x"81ff0bd4",
   248 => x"0c81ff0b",
   249 => x"d40c81ff",
   250 => x"0bd40c72",
   251 => x"862a7081",
   252 => x"06a4c008",
   253 => x"56515372",
   254 => x"802eff84",
   255 => x"38810ba4",
   256 => x"c00c0290",
   257 => x"050d0402",
   258 => x"e8050d78",
   259 => x"5681ff0b",
   260 => x"d40cd008",
   261 => x"708f2a70",
   262 => x"81065151",
   263 => x"5372f338",
   264 => x"82810bd0",
   265 => x"0c81ff0b",
   266 => x"d40c7752",
   267 => x"87fc80d8",
   268 => x"5184b42d",
   269 => x"a4c00881",
   270 => x"823881ff",
   271 => x"0bd40c81",
   272 => x"fe0bd40c",
   273 => x"80ff5575",
   274 => x"70840557",
   275 => x"0870982a",
   276 => x"d40c7090",
   277 => x"2c7081ff",
   278 => x"06d40c54",
   279 => x"70882c70",
   280 => x"81ff06d4",
   281 => x"0c547081",
   282 => x"ff06d40c",
   283 => x"54ff1555",
   284 => x"748025d3",
   285 => x"3881ff0b",
   286 => x"d40c81ff",
   287 => x"0bd40c81",
   288 => x"ff0bd40c",
   289 => x"868da054",
   290 => x"81ff0bd4",
   291 => x"0cd40881",
   292 => x"ff065574",
   293 => x"8738ff14",
   294 => x"5473ed38",
   295 => x"81ff0bd4",
   296 => x"0cd00870",
   297 => x"8f2a7081",
   298 => x"06515153",
   299 => x"72f33872",
   300 => x"d00c72a4",
   301 => x"c00c0298",
   302 => x"050d04a2",
   303 => x"c851839e",
   304 => x"2d810ba4",
   305 => x"c00c0298",
   306 => x"050d0402",
   307 => x"ec050d76",
   308 => x"78545480",
   309 => x"5580dbc6",
   310 => x"df5281ff",
   311 => x"0bd40cd4",
   312 => x"087081ff",
   313 => x"06515170",
   314 => x"81fe2e95",
   315 => x"38ff1252",
   316 => x"71e83881",
   317 => x"ff0bd40c",
   318 => x"74a4c00c",
   319 => x"0294050d",
   320 => x"04800ba5",
   321 => x"c80c8373",
   322 => x"259f3883",
   323 => x"e62da4c0",
   324 => x"08747084",
   325 => x"05560ca5",
   326 => x"c808a4c0",
   327 => x"0805a5c8",
   328 => x"0cfc1353",
   329 => x"728324e3",
   330 => x"38807325",
   331 => x"a03881ff",
   332 => x"0bd40cff",
   333 => x"74708105",
   334 => x"5681b72d",
   335 => x"a5c80881",
   336 => x"ff05a5c8",
   337 => x"0cff1353",
   338 => x"728024e2",
   339 => x"38815581",
   340 => x"ff0bd40c",
   341 => x"74a4c00c",
   342 => x"0294050d",
   343 => x"0402e805",
   344 => x"0d805287",
   345 => x"fc80c951",
   346 => x"84b42d92",
   347 => x"52a5b451",
   348 => x"89cb2da5",
   349 => x"b40b80f5",
   350 => x"2d81c006",
   351 => x"537280c0",
   352 => x"2e80f738",
   353 => x"a5bd0b80",
   354 => x"f52d7010",
   355 => x"8606a5be",
   356 => x"0b80f52d",
   357 => x"70872a72",
   358 => x"07a5b90b",
   359 => x"80f52d8f",
   360 => x"06a5ba0b",
   361 => x"80f52d70",
   362 => x"8a2b9880",
   363 => x"06a5bb0b",
   364 => x"80f52d70",
   365 => x"822b7207",
   366 => x"a5bc0b80",
   367 => x"f52d7086",
   368 => x"2a720782",
   369 => x"1881782b",
   370 => x"81138173",
   371 => x"2b712951",
   372 => x"53585852",
   373 => x"52525259",
   374 => x"53545258",
   375 => x"55558480",
   376 => x"75258e38",
   377 => x"72107581",
   378 => x"2c565374",
   379 => x"848024f4",
   380 => x"3872a4c0",
   381 => x"0c029805",
   382 => x"0d04a5bb",
   383 => x"0b80f52d",
   384 => x"a5bc0b80",
   385 => x"f52d7190",
   386 => x"2b71882b",
   387 => x"07a5bd0b",
   388 => x"80f52d71",
   389 => x"81fffe80",
   390 => x"06077088",
   391 => x"80298880",
   392 => x"05a4c00c",
   393 => x"51555755",
   394 => x"0298050d",
   395 => x"0402f005",
   396 => x"0d810ba5",
   397 => x"a40ca2d8",
   398 => x"51839e2d",
   399 => x"8754d008",
   400 => x"708f2a70",
   401 => x"81065151",
   402 => x"5372f338",
   403 => x"72d00c85",
   404 => x"a52dd008",
   405 => x"708f2a70",
   406 => x"81065151",
   407 => x"5372f338",
   408 => x"810bd00c",
   409 => x"725284d4",
   410 => x"80c05184",
   411 => x"b42da4c0",
   412 => x"08812e8e",
   413 => x"3873822e",
   414 => x"80e138ff",
   415 => x"145473ff",
   416 => x"bd3886e2",
   417 => x"2da4c008",
   418 => x"a5a40ca4",
   419 => x"c008802e",
   420 => x"af3881ff",
   421 => x"0bd40c8a",
   422 => x"dd2da4c0",
   423 => x"08a5a80c",
   424 => x"d008708f",
   425 => x"2a708106",
   426 => x"51515372",
   427 => x"f33872d0",
   428 => x"0c81ff0b",
   429 => x"d40c810b",
   430 => x"a4c00c02",
   431 => x"90050d04",
   432 => x"815287fc",
   433 => x"80d05184",
   434 => x"b42d81ff",
   435 => x"0bd40c8a",
   436 => x"dd2da4c0",
   437 => x"08a5a80c",
   438 => x"8da004a2",
   439 => x"dc51839e",
   440 => x"2d72a4c0",
   441 => x"0c029005",
   442 => x"0d0402f0",
   443 => x"050d8054",
   444 => x"81ff0bd4",
   445 => x"0cd00870",
   446 => x"8f2a7081",
   447 => x"06515153",
   448 => x"72f33882",
   449 => x"810bd00c",
   450 => x"81ff0bd4",
   451 => x"0c755287",
   452 => x"fc80d151",
   453 => x"84b42da4",
   454 => x"c008802e",
   455 => x"8a3873a4",
   456 => x"c00c0290",
   457 => x"050d0484",
   458 => x"80527651",
   459 => x"89cb2da4",
   460 => x"c00854d0",
   461 => x"08708f2a",
   462 => x"70810651",
   463 => x"515372f3",
   464 => x"3872d00c",
   465 => x"73a4c00c",
   466 => x"0290050d",
   467 => x"0402f405",
   468 => x"0d747088",
   469 => x"2a83fe80",
   470 => x"06707298",
   471 => x"2a077288",
   472 => x"2b87fc80",
   473 => x"80067398",
   474 => x"2b81f00a",
   475 => x"06717307",
   476 => x"07a4c00c",
   477 => x"56515351",
   478 => x"028c050d",
   479 => x"0402f805",
   480 => x"0d028e05",
   481 => x"80f52d74",
   482 => x"882b0770",
   483 => x"83ffff06",
   484 => x"a4c00c51",
   485 => x"0288050d",
   486 => x"0402f805",
   487 => x"0d737090",
   488 => x"2b71902a",
   489 => x"07a4c00c",
   490 => x"52028805",
   491 => x"0d0402f4",
   492 => x"050da5a0",
   493 => x"0853cc08",
   494 => x"70828006",
   495 => x"52527073",
   496 => x"2ef43872",
   497 => x"828032a5",
   498 => x"a00c71fd",
   499 => x"ff06a4c0",
   500 => x"0c028c05",
   501 => x"0d0402d8",
   502 => x"050d800b",
   503 => x"a5a00ca2",
   504 => x"e451839e",
   505 => x"2d8cad2d",
   506 => x"a4c0088b",
   507 => x"38800ba4",
   508 => x"c00c02a8",
   509 => x"050d04a2",
   510 => x"ec51839e",
   511 => x"2d96eb2d",
   512 => x"8fae2da4",
   513 => x"c0085aa4",
   514 => x"c0088182",
   515 => x"2e80c438",
   516 => x"a4c00881",
   517 => x"822482ec",
   518 => x"38a4c008",
   519 => x"842e83a8",
   520 => x"38a4c008",
   521 => x"842484e1",
   522 => x"38a4c008",
   523 => x"832e80e5",
   524 => x"38905380",
   525 => x"52795181",
   526 => x"f72da2f4",
   527 => x"51839e2d",
   528 => x"8fae2da4",
   529 => x"c0085aa4",
   530 => x"c0088182",
   531 => x"2e098106",
   532 => x"ffbe38a2",
   533 => x"f851839e",
   534 => x"2da5a80b",
   535 => x"80f52da5",
   536 => x"a00807cc",
   537 => x"0c8fae2d",
   538 => x"a5a90b80",
   539 => x"f52da5a0",
   540 => x"0807cc0c",
   541 => x"8fae2da5",
   542 => x"aa0b80f5",
   543 => x"2da5a008",
   544 => x"07cc0c8f",
   545 => x"ae2da5ab",
   546 => x"0b80f52d",
   547 => x"a5a00807",
   548 => x"cc0c9080",
   549 => x"0480f251",
   550 => x"82da2da5",
   551 => x"a008cc0c",
   552 => x"8fae2da4",
   553 => x"c008982b",
   554 => x"a5a008cc",
   555 => x"0c588fae",
   556 => x"2da4c008",
   557 => x"902b7807",
   558 => x"a5a008cc",
   559 => x"0c588fae",
   560 => x"2da4c008",
   561 => x"882b7807",
   562 => x"a5a008cc",
   563 => x"0c588fae",
   564 => x"2d77a4c0",
   565 => x"0807a5a0",
   566 => x"08cc0c58",
   567 => x"8fae2da4",
   568 => x"c008ff05",
   569 => x"5978ff2e",
   570 => x"80f438a5",
   571 => x"e4577983",
   572 => x"2e80f338",
   573 => x"76527751",
   574 => x"8118588d",
   575 => x"ea2d80ff",
   576 => x"56767084",
   577 => x"05580870",
   578 => x"982aa5a0",
   579 => x"0807cc0c",
   580 => x"558fae2d",
   581 => x"74902a70",
   582 => x"81ff0670",
   583 => x"a5a00807",
   584 => x"cc0c5154",
   585 => x"8fae2d74",
   586 => x"882a7081",
   587 => x"ff0670a5",
   588 => x"a00807cc",
   589 => x"0c51548f",
   590 => x"ae2d7481",
   591 => x"ff0670a5",
   592 => x"a00807cc",
   593 => x"0c558fae",
   594 => x"2dff1656",
   595 => x"758025ff",
   596 => x"b038ff19",
   597 => x"5978ff2e",
   598 => x"098106ff",
   599 => x"8e38a5a0",
   600 => x"08cc0c90",
   601 => x"8004a051",
   602 => x"82da2d77",
   603 => x"528118a9",
   604 => x"e85258a0",
   605 => x"ff2d7652",
   606 => x"a9e851a0",
   607 => x"912d80ff",
   608 => x"56928104",
   609 => x"a4c00881",
   610 => x"842ebd38",
   611 => x"81840ba4",
   612 => x"c00824fe",
   613 => x"8038a4c0",
   614 => x"0881902e",
   615 => x"828238a4",
   616 => x"c00881fe",
   617 => x"2e098106",
   618 => x"fd8738a5",
   619 => x"a00881fe",
   620 => x"07cc0c8f",
   621 => x"ae2da4c0",
   622 => x"085182da",
   623 => x"2da5a008",
   624 => x"81fe07cc",
   625 => x"0c908004",
   626 => x"a5a008cc",
   627 => x"0c8fae2d",
   628 => x"a4c00898",
   629 => x"2ba5a008",
   630 => x"cc0c588f",
   631 => x"ae2da4c0",
   632 => x"08902b78",
   633 => x"07a5a008",
   634 => x"cc0c588f",
   635 => x"ae2da4c0",
   636 => x"08882b78",
   637 => x"07a5a008",
   638 => x"cc0c588f",
   639 => x"ae2d77a4",
   640 => x"c00807a5",
   641 => x"a008cc0c",
   642 => x"588fae2d",
   643 => x"a4c00859",
   644 => x"80f75182",
   645 => x"da2dff19",
   646 => x"5978ff2e",
   647 => x"fec038a5",
   648 => x"e4557984",
   649 => x"2e81c438",
   650 => x"80ff56a5",
   651 => x"a008cc0c",
   652 => x"8fae2da5",
   653 => x"a008cc0c",
   654 => x"a4c00888",
   655 => x"2b548fae",
   656 => x"2da5a008",
   657 => x"cc0c73a4",
   658 => x"c0080788",
   659 => x"2b548fae",
   660 => x"2da5a008",
   661 => x"cc0c73a4",
   662 => x"c0080788",
   663 => x"2b548fae",
   664 => x"2d73a4c0",
   665 => x"08077570",
   666 => x"8405570c",
   667 => x"ff165675",
   668 => x"8025ffb7",
   669 => x"3879842e",
   670 => x"818238a5",
   671 => x"e4527751",
   672 => x"81185888",
   673 => x"872d9496",
   674 => x"04a4c008",
   675 => x"81802e09",
   676 => x"8106fb9d",
   677 => x"38a5a008",
   678 => x"818007cc",
   679 => x"0c908004",
   680 => x"8056a5a0",
   681 => x"08cc0ca5",
   682 => x"cc16548f",
   683 => x"ae2da4c0",
   684 => x"087481b7",
   685 => x"2d811656",
   686 => x"8b7625e6",
   687 => x"38800ba5",
   688 => x"d70b81b7",
   689 => x"2da5cc51",
   690 => x"839e2da5",
   691 => x"cc52a9e8",
   692 => x"519d9a2d",
   693 => x"a4c00880",
   694 => x"2eae38a5",
   695 => x"a008cc0c",
   696 => x"8fae2da5",
   697 => x"a008cc0c",
   698 => x"90800477",
   699 => x"528118a9",
   700 => x"e85258a0",
   701 => x"ff2d80ff",
   702 => x"5694ab04",
   703 => x"a5e452a9",
   704 => x"e851a0c8",
   705 => x"2d949604",
   706 => x"a5a00881",
   707 => x"ff07cc0c",
   708 => x"8fae2da5",
   709 => x"a00881ff",
   710 => x"07cc0ca3",
   711 => x"8051839e",
   712 => x"2d90c004",
   713 => x"02e8050d",
   714 => x"77797b58",
   715 => x"55558053",
   716 => x"727625a3",
   717 => x"38747081",
   718 => x"055680f5",
   719 => x"2d747081",
   720 => x"055680f5",
   721 => x"2d525271",
   722 => x"712e0981",
   723 => x"06933881",
   724 => x"13537573",
   725 => x"24df3880",
   726 => x"0ba4c00c",
   727 => x"0298050d",
   728 => x"04810ba4",
   729 => x"c00c0298",
   730 => x"050d0402",
   731 => x"d8050d80",
   732 => x"0baa8c0c",
   733 => x"a3885183",
   734 => x"9e2da5e4",
   735 => x"5280518d",
   736 => x"ea2da4c0",
   737 => x"0854a4c0",
   738 => x"089238a3",
   739 => x"9851839e",
   740 => x"2d735675",
   741 => x"a4c00c02",
   742 => x"a8050d04",
   743 => x"a3ac5183",
   744 => x"9e2d8055",
   745 => x"810ba5d8",
   746 => x"0c8853a3",
   747 => x"c452a69a",
   748 => x"5196a42d",
   749 => x"a4c00875",
   750 => x"2e80fb38",
   751 => x"8853a3d0",
   752 => x"52a6b651",
   753 => x"96a42da4",
   754 => x"c0088738",
   755 => x"a4c008a5",
   756 => x"d80ca5d8",
   757 => x"08802e81",
   758 => x"8938a9aa",
   759 => x"0b80f52d",
   760 => x"a9ab0b80",
   761 => x"f52d7198",
   762 => x"2b71902b",
   763 => x"07a9ac0b",
   764 => x"80f52d70",
   765 => x"882b7207",
   766 => x"a9ad0b80",
   767 => x"f52d7107",
   768 => x"a9e20b80",
   769 => x"f52da9e3",
   770 => x"0b80f52d",
   771 => x"71882b07",
   772 => x"53405552",
   773 => x"5a565755",
   774 => x"7381abaa",
   775 => x"2ea13873",
   776 => x"82d4d52e",
   777 => x"a338a3dc",
   778 => x"51839e2d",
   779 => x"800ba4c0",
   780 => x"0c02a805",
   781 => x"0d04a4c0",
   782 => x"08a5d80c",
   783 => x"97bc0474",
   784 => x"518ecd2d",
   785 => x"a4c00855",
   786 => x"a5e45274",
   787 => x"518dea2d",
   788 => x"a4c00856",
   789 => x"a4c00880",
   790 => x"2efeb838",
   791 => x"a3fc5183",
   792 => x"9e2d8853",
   793 => x"a3d052a6",
   794 => x"b65196a4",
   795 => x"2da4c008",
   796 => x"81fa3881",
   797 => x"0baa8c0c",
   798 => x"a9e20b80",
   799 => x"f52d5473",
   800 => x"80d52e09",
   801 => x"8106ffa4",
   802 => x"38a9e30b",
   803 => x"80f52d54",
   804 => x"7381aa2e",
   805 => x"098106ff",
   806 => x"9338800b",
   807 => x"a5e40b80",
   808 => x"f52d5754",
   809 => x"7581e92e",
   810 => x"83388154",
   811 => x"7581eb2e",
   812 => x"8c388056",
   813 => x"73762e09",
   814 => x"8106fdd7",
   815 => x"38a5ef0b",
   816 => x"80f52d56",
   817 => x"75fee538",
   818 => x"a5f00b80",
   819 => x"f52d5473",
   820 => x"822e0981",
   821 => x"06fed538",
   822 => x"a5f10b80",
   823 => x"f52d70aa",
   824 => x"940cff05",
   825 => x"aa880ca5",
   826 => x"f20b80f5",
   827 => x"2da5f30b",
   828 => x"80f52d5b",
   829 => x"75057a82",
   830 => x"80290570",
   831 => x"a9fc0ca5",
   832 => x"f40b80f5",
   833 => x"2d70a9f8",
   834 => x"0caa8c08",
   835 => x"5b595778",
   836 => x"80f838a5",
   837 => x"f60b80f5",
   838 => x"2da5f50b",
   839 => x"80f52d71",
   840 => x"82802905",
   841 => x"70a9e40c",
   842 => x"70a02983",
   843 => x"ff057089",
   844 => x"2a70aa90",
   845 => x"0ca5fb0b",
   846 => x"80f52da5",
   847 => x"fa0b80f5",
   848 => x"2d718280",
   849 => x"290570a5",
   850 => x"dc0c7d71",
   851 => x"291d70aa",
   852 => x"840c7fa5",
   853 => x"e00c7305",
   854 => x"aa9c0c5a",
   855 => x"5a515155",
   856 => x"5a815675",
   857 => x"a4c00c02",
   858 => x"a8050d04",
   859 => x"8853a3c4",
   860 => x"52a69a51",
   861 => x"96a42d80",
   862 => x"56a4c008",
   863 => x"762efdf8",
   864 => x"3875a4c0",
   865 => x"0c02a805",
   866 => x"0d048853",
   867 => x"a3d052a6",
   868 => x"b65196a4",
   869 => x"2da4c008",
   870 => x"fbf938aa",
   871 => x"94087084",
   872 => x"2ba9e40c",
   873 => x"70aa900c",
   874 => x"a6890b80",
   875 => x"f52da688",
   876 => x"0b80f52d",
   877 => x"71828029",
   878 => x"05a68a0b",
   879 => x"80f52d70",
   880 => x"84808029",
   881 => x"12a68b0b",
   882 => x"80f52d70",
   883 => x"81800a29",
   884 => x"1270a5dc",
   885 => x"0ca9f808",
   886 => x"7129a9fc",
   887 => x"080570aa",
   888 => x"9c0ca691",
   889 => x"0b80f52d",
   890 => x"a6900b80",
   891 => x"f52d7182",
   892 => x"802905a6",
   893 => x"920b80f5",
   894 => x"2d708480",
   895 => x"802912a6",
   896 => x"930b80f5",
   897 => x"2d70982b",
   898 => x"81f00a06",
   899 => x"720570a5",
   900 => x"e00cfe11",
   901 => x"7e297705",
   902 => x"aa840c52",
   903 => x"59525558",
   904 => x"5e51525f",
   905 => x"525b5755",
   906 => x"5781569a",
   907 => x"e30402ec",
   908 => x"050d7670",
   909 => x"872c7180",
   910 => x"ff065656",
   911 => x"53aa8c08",
   912 => x"8a387288",
   913 => x"2c7381ff",
   914 => x"065555a5",
   915 => x"e452a9fc",
   916 => x"0815518d",
   917 => x"ea2da4c0",
   918 => x"0853a4c0",
   919 => x"08802e9c",
   920 => x"38aa8c08",
   921 => x"802e9e38",
   922 => x"731010a5",
   923 => x"e4057008",
   924 => x"52538ecd",
   925 => x"2da4c008",
   926 => x"f00a0653",
   927 => x"72a4c00c",
   928 => x"0294050d",
   929 => x"047310a5",
   930 => x"e4057080",
   931 => x"e02d5253",
   932 => x"8efd2da4",
   933 => x"c008539c",
   934 => x"fc0402cc",
   935 => x"050d7e60",
   936 => x"5d5d800b",
   937 => x"a5e008aa",
   938 => x"84085a5c",
   939 => x"57aa8c08",
   940 => x"772e818a",
   941 => x"38aa9408",
   942 => x"842b5980",
   943 => x"56757927",
   944 => x"80c43875",
   945 => x"8f06a018",
   946 => x"58547380",
   947 => x"2e80fa38",
   948 => x"807780f5",
   949 => x"2d555573",
   950 => x"752e8338",
   951 => x"81557381",
   952 => x"e52e9a38",
   953 => x"81707606",
   954 => x"555a7380",
   955 => x"2e8f388b",
   956 => x"1780f52d",
   957 => x"98065574",
   958 => x"802e80de",
   959 => x"38811656",
   960 => x"787626ff",
   961 => x"be38aa8c",
   962 => x"08802e81",
   963 => x"c1387a51",
   964 => x"9cae2da4",
   965 => x"c008a4c0",
   966 => x"0880ffff",
   967 => x"fff80655",
   968 => x"5b7380ff",
   969 => x"fffff82e",
   970 => x"81a438a4",
   971 => x"c008fe05",
   972 => x"aa940829",
   973 => x"aa9c0805",
   974 => x"5880569d",
   975 => x"bd04aa90",
   976 => x"08842b59",
   977 => x"80569dbd",
   978 => x"04a5e452",
   979 => x"77518118",
   980 => x"588dea2d",
   981 => x"a5e4579d",
   982 => x"d0048b53",
   983 => x"7b527651",
   984 => x"96a42da4",
   985 => x"c008ff95",
   986 => x"389c1708",
   987 => x"518ecd2d",
   988 => x"a4c00884",
   989 => x"1e0c9a17",
   990 => x"80e02d51",
   991 => x"8efd2da4",
   992 => x"c008a4c0",
   993 => x"085556aa",
   994 => x"8c089738",
   995 => x"73881e0c",
   996 => x"738c1e0c",
   997 => x"747d0c79",
   998 => x"5473a4c0",
   999 => x"0c02b405",
  1000 => x"0d04a4c0",
  1001 => x"08881e0c",
  1002 => x"941780e0",
  1003 => x"2d518efd",
  1004 => x"2da4c008",
  1005 => x"902b83ff",
  1006 => x"f00a0670",
  1007 => x"17707f88",
  1008 => x"050c8c1f",
  1009 => x"0c54747d",
  1010 => x"0c79549f",
  1011 => x"9904800b",
  1012 => x"a4c00c02",
  1013 => x"b4050d04",
  1014 => x"02f4050d",
  1015 => x"74700881",
  1016 => x"05710c70",
  1017 => x"08aa8808",
  1018 => x"06535371",
  1019 => x"802e8b38",
  1020 => x"810ba4c0",
  1021 => x"0c028c05",
  1022 => x"0d048813",
  1023 => x"08519cae",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


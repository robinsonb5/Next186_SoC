-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba4",
     9 => x"b0080b0b",
    10 => x"0ba4b408",
    11 => x"0b0b0ba4",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a4b80c0b",
    16 => x"0b0ba4b4",
    17 => x"0c0b0b0b",
    18 => x"a4b00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba2ac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a4b070aa",
    57 => x"90278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8fd00402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752e80c7",
    65 => x"38875472",
    66 => x"9c2a7384",
    67 => x"2b545271",
    68 => x"802e8338",
    69 => x"81558972",
    70 => x"259938b7",
    71 => x"1252749b",
    72 => x"38ff1454",
    73 => x"738025df",
    74 => x"38800ba4",
    75 => x"b00c0294",
    76 => x"050d04b0",
    77 => x"12527480",
    78 => x"2ee73871",
    79 => x"5182da2d",
    80 => x"ff145473",
    81 => x"8025c038",
    82 => x"82a904b0",
    83 => x"5182da2d",
    84 => x"800ba4b0",
    85 => x"0c029405",
    86 => x"0d0402f8",
    87 => x"050d7352",
    88 => x"c0087088",
    89 => x"2a708106",
    90 => x"51515170",
    91 => x"802ef138",
    92 => x"71c00c71",
    93 => x"a4b00c02",
    94 => x"88050d04",
    95 => x"02f8050d",
    96 => x"7352c408",
    97 => x"70882a70",
    98 => x"81065151",
    99 => x"5170802e",
   100 => x"f13871c4",
   101 => x"0c71a4b0",
   102 => x"0c028805",
   103 => x"0d0402e8",
   104 => x"050d8078",
   105 => x"57557570",
   106 => x"84055708",
   107 => x"53805472",
   108 => x"982a7388",
   109 => x"2b545271",
   110 => x"802ea238",
   111 => x"c0087088",
   112 => x"2a708106",
   113 => x"51515170",
   114 => x"802ef138",
   115 => x"71c00c81",
   116 => x"15811555",
   117 => x"55837425",
   118 => x"d63871ca",
   119 => x"3874a4b0",
   120 => x"0c029805",
   121 => x"0d0402f4",
   122 => x"050dd452",
   123 => x"81ff720c",
   124 => x"71085381",
   125 => x"ff720c72",
   126 => x"882b83fe",
   127 => x"80067208",
   128 => x"7081ff06",
   129 => x"51525381",
   130 => x"ff720c72",
   131 => x"7107882b",
   132 => x"72087081",
   133 => x"ff065152",
   134 => x"5381ff72",
   135 => x"0c727107",
   136 => x"882b7208",
   137 => x"7081ff06",
   138 => x"7207a4b0",
   139 => x"0c525302",
   140 => x"8c050d04",
   141 => x"02f4050d",
   142 => x"74767181",
   143 => x"ff06d40c",
   144 => x"5353a594",
   145 => x"08853871",
   146 => x"892b5271",
   147 => x"982ad40c",
   148 => x"71902a70",
   149 => x"81ff06d4",
   150 => x"0c517188",
   151 => x"2a7081ff",
   152 => x"06d40c51",
   153 => x"7181ff06",
   154 => x"d40c7290",
   155 => x"2a7081ff",
   156 => x"06d40c51",
   157 => x"d4087081",
   158 => x"ff065151",
   159 => x"82b8bf52",
   160 => x"7081ff2e",
   161 => x"09810694",
   162 => x"3881ff0b",
   163 => x"d40cd408",
   164 => x"7081ff06",
   165 => x"ff145451",
   166 => x"5171e538",
   167 => x"70a4b00c",
   168 => x"028c050d",
   169 => x"0402fc05",
   170 => x"0d81c751",
   171 => x"81ff0bd4",
   172 => x"0cff1151",
   173 => x"708025f4",
   174 => x"38028405",
   175 => x"0d0402f0",
   176 => x"050d85a5",
   177 => x"2d819c9f",
   178 => x"53805287",
   179 => x"fc80f751",
   180 => x"84b42da4",
   181 => x"b00854a4",
   182 => x"b008812e",
   183 => x"9038ff13",
   184 => x"5372e638",
   185 => x"72a4b00c",
   186 => x"0290050d",
   187 => x"0481ff0b",
   188 => x"d40c820a",
   189 => x"52849c80",
   190 => x"e95184b4",
   191 => x"2da4b008",
   192 => x"802e8e38",
   193 => x"85a52dff",
   194 => x"135372ff",
   195 => x"bc3885e4",
   196 => x"0481ff0b",
   197 => x"d40c73a4",
   198 => x"b00c0290",
   199 => x"050d0402",
   200 => x"f4050d81",
   201 => x"ff0bd40c",
   202 => x"a2bc5183",
   203 => x"9e2d9353",
   204 => x"805287fc",
   205 => x"80c15184",
   206 => x"b42da4b0",
   207 => x"08802e93",
   208 => x"3885a52d",
   209 => x"ff135372",
   210 => x"e73872a4",
   211 => x"b00c028c",
   212 => x"050d0481",
   213 => x"ff0bd40c",
   214 => x"810ba4b0",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050d85a5",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"5184b42d",
   221 => x"a4b00881",
   222 => x"2e8f3886",
   223 => x"9f2d8054",
   224 => x"73a4b00c",
   225 => x"0290050d",
   226 => x"0483e62d",
   227 => x"a4b00883",
   228 => x"ffff0653",
   229 => x"7283aa2e",
   230 => x"098106df",
   231 => x"3881ff0b",
   232 => x"d40cb153",
   233 => x"85be2da4",
   234 => x"b0089538",
   235 => x"72822ece",
   236 => x"38ff1353",
   237 => x"72ee3872",
   238 => x"a4b00c02",
   239 => x"90050d04",
   240 => x"805287fc",
   241 => x"80fa5184",
   242 => x"b42da4b0",
   243 => x"08de3881",
   244 => x"ff0bd40c",
   245 => x"d4085381",
   246 => x"ff0bd40c",
   247 => x"81ff0bd4",
   248 => x"0c81ff0b",
   249 => x"d40c81ff",
   250 => x"0bd40c72",
   251 => x"862a7081",
   252 => x"06a4b008",
   253 => x"56515372",
   254 => x"802eff84",
   255 => x"38810ba4",
   256 => x"b00c0290",
   257 => x"050d0402",
   258 => x"e8050d78",
   259 => x"5681ff0b",
   260 => x"d40cd008",
   261 => x"708f2a70",
   262 => x"81065151",
   263 => x"5372f338",
   264 => x"82810bd0",
   265 => x"0c81ff0b",
   266 => x"d40c7752",
   267 => x"87fc80d8",
   268 => x"5184b42d",
   269 => x"a4b00881",
   270 => x"823881ff",
   271 => x"0bd40c81",
   272 => x"fe0bd40c",
   273 => x"80ff5575",
   274 => x"70840557",
   275 => x"0870982a",
   276 => x"d40c7090",
   277 => x"2c7081ff",
   278 => x"06d40c54",
   279 => x"70882c70",
   280 => x"81ff06d4",
   281 => x"0c547081",
   282 => x"ff06d40c",
   283 => x"54ff1555",
   284 => x"748025d3",
   285 => x"3881ff0b",
   286 => x"d40c81ff",
   287 => x"0bd40c81",
   288 => x"ff0bd40c",
   289 => x"868da054",
   290 => x"81ff0bd4",
   291 => x"0cd40881",
   292 => x"ff065574",
   293 => x"8738ff14",
   294 => x"5473ed38",
   295 => x"81ff0bd4",
   296 => x"0cd00870",
   297 => x"8f2a7081",
   298 => x"06515153",
   299 => x"72f33872",
   300 => x"d00c72a4",
   301 => x"b00c0298",
   302 => x"050d04a2",
   303 => x"c051839e",
   304 => x"2d810ba4",
   305 => x"b00c0298",
   306 => x"050d0402",
   307 => x"ec050d76",
   308 => x"78545480",
   309 => x"5580dbc6",
   310 => x"df5281ff",
   311 => x"0bd40cd4",
   312 => x"087081ff",
   313 => x"06515170",
   314 => x"81fe2e95",
   315 => x"38ff1252",
   316 => x"71e83881",
   317 => x"ff0bd40c",
   318 => x"74a4b00c",
   319 => x"0294050d",
   320 => x"04800ba5",
   321 => x"b80c8373",
   322 => x"259f3883",
   323 => x"e62da4b0",
   324 => x"08747084",
   325 => x"05560ca5",
   326 => x"b808a4b0",
   327 => x"0805a5b8",
   328 => x"0cfc1353",
   329 => x"728324e3",
   330 => x"38807325",
   331 => x"a03881ff",
   332 => x"0bd40cff",
   333 => x"74708105",
   334 => x"5681b72d",
   335 => x"a5b80881",
   336 => x"ff05a5b8",
   337 => x"0cff1353",
   338 => x"728024e2",
   339 => x"38815581",
   340 => x"ff0bd40c",
   341 => x"74a4b00c",
   342 => x"0294050d",
   343 => x"0402e805",
   344 => x"0d805287",
   345 => x"fc80c951",
   346 => x"84b42d92",
   347 => x"52a5a451",
   348 => x"89cb2da5",
   349 => x"a40b80f5",
   350 => x"2d81c006",
   351 => x"537280c0",
   352 => x"2e80f738",
   353 => x"a5ad0b80",
   354 => x"f52d7010",
   355 => x"8606a5ae",
   356 => x"0b80f52d",
   357 => x"70872a72",
   358 => x"07a5a90b",
   359 => x"80f52d8f",
   360 => x"06a5aa0b",
   361 => x"80f52d70",
   362 => x"8a2b9880",
   363 => x"06a5ab0b",
   364 => x"80f52d70",
   365 => x"822b7207",
   366 => x"a5ac0b80",
   367 => x"f52d7086",
   368 => x"2a720782",
   369 => x"1881782b",
   370 => x"81138173",
   371 => x"2b712951",
   372 => x"53585852",
   373 => x"52525259",
   374 => x"53545258",
   375 => x"55558480",
   376 => x"75258e38",
   377 => x"72107581",
   378 => x"2c565374",
   379 => x"848024f4",
   380 => x"3872a4b0",
   381 => x"0c029805",
   382 => x"0d04a5ab",
   383 => x"0b80f52d",
   384 => x"a5ac0b80",
   385 => x"f52d7190",
   386 => x"2b71882b",
   387 => x"07a5ad0b",
   388 => x"80f52d71",
   389 => x"81fffe80",
   390 => x"06077088",
   391 => x"80298880",
   392 => x"05a4b00c",
   393 => x"51555755",
   394 => x"0298050d",
   395 => x"0402f405",
   396 => x"0d810ba5",
   397 => x"940cd008",
   398 => x"708f2a70",
   399 => x"81065151",
   400 => x"5372f338",
   401 => x"72d00c85",
   402 => x"a52da2d0",
   403 => x"51839e2d",
   404 => x"d008708f",
   405 => x"2a708106",
   406 => x"51515372",
   407 => x"f338810b",
   408 => x"d00c8753",
   409 => x"805284d4",
   410 => x"80c05184",
   411 => x"b42da4b0",
   412 => x"08812e8d",
   413 => x"3872822e",
   414 => x"80c538ff",
   415 => x"135372e4",
   416 => x"3886e22d",
   417 => x"a4b008a5",
   418 => x"940ca4b0",
   419 => x"08802eb9",
   420 => x"3881ff0b",
   421 => x"d40c8add",
   422 => x"2da4b008",
   423 => x"a5980cd0",
   424 => x"08708f2a",
   425 => x"70810651",
   426 => x"515372f3",
   427 => x"3872d00c",
   428 => x"81ff0bd4",
   429 => x"0c810ba4",
   430 => x"b00c028c",
   431 => x"050d0480",
   432 => x"0ba4b00c",
   433 => x"028c050d",
   434 => x"04815287",
   435 => x"fc80d051",
   436 => x"84b42d81",
   437 => x"ff0bd40c",
   438 => x"8add2da4",
   439 => x"b008a598",
   440 => x"0c8d9f04",
   441 => x"02f0050d",
   442 => x"805481ff",
   443 => x"0bd40cd0",
   444 => x"08708f2a",
   445 => x"70810651",
   446 => x"515372f3",
   447 => x"3882810b",
   448 => x"d00c81ff",
   449 => x"0bd40c75",
   450 => x"5287fc80",
   451 => x"d15184b4",
   452 => x"2da4b008",
   453 => x"802e8a38",
   454 => x"73a4b00c",
   455 => x"0290050d",
   456 => x"04848052",
   457 => x"765189cb",
   458 => x"2da4b008",
   459 => x"54d00870",
   460 => x"8f2a7081",
   461 => x"06515153",
   462 => x"72f33872",
   463 => x"d00c73a4",
   464 => x"b00c0290",
   465 => x"050d0402",
   466 => x"f4050d74",
   467 => x"70882a83",
   468 => x"fe800670",
   469 => x"72982a07",
   470 => x"72882b87",
   471 => x"fc808006",
   472 => x"73982b81",
   473 => x"f00a0671",
   474 => x"730707a4",
   475 => x"b00c5651",
   476 => x"5351028c",
   477 => x"050d0402",
   478 => x"f8050d02",
   479 => x"8e0580f5",
   480 => x"2d74882b",
   481 => x"077083ff",
   482 => x"ff06a4b0",
   483 => x"0c510288",
   484 => x"050d0402",
   485 => x"f8050d73",
   486 => x"70902b71",
   487 => x"902a07a4",
   488 => x"b00c5202",
   489 => x"88050d04",
   490 => x"02f4050d",
   491 => x"a5900853",
   492 => x"cc087082",
   493 => x"80065252",
   494 => x"70732ef4",
   495 => x"38728280",
   496 => x"32a5900c",
   497 => x"71fdff06",
   498 => x"a4b00c02",
   499 => x"8c050d04",
   500 => x"02d8050d",
   501 => x"800ba590",
   502 => x"0ca2d451",
   503 => x"839e2d8c",
   504 => x"ad2da4b0",
   505 => x"088b3880",
   506 => x"0ba4b00c",
   507 => x"02a8050d",
   508 => x"04a2dc51",
   509 => x"839e2d96",
   510 => x"e52d8fa8",
   511 => x"2da4b008",
   512 => x"5aa4b008",
   513 => x"81822e80",
   514 => x"c438a4b0",
   515 => x"08818224",
   516 => x"82ec38a4",
   517 => x"b008842e",
   518 => x"83a838a4",
   519 => x"b0088424",
   520 => x"84e138a4",
   521 => x"b008832e",
   522 => x"80e53890",
   523 => x"53805279",
   524 => x"5181f72d",
   525 => x"a2e45183",
   526 => x"9e2d8fa8",
   527 => x"2da4b008",
   528 => x"5aa4b008",
   529 => x"81822e09",
   530 => x"8106ffbe",
   531 => x"38a2e851",
   532 => x"839e2da5",
   533 => x"980b80f5",
   534 => x"2da59008",
   535 => x"07cc0c8f",
   536 => x"a82da599",
   537 => x"0b80f52d",
   538 => x"a5900807",
   539 => x"cc0c8fa8",
   540 => x"2da59a0b",
   541 => x"80f52da5",
   542 => x"900807cc",
   543 => x"0c8fa82d",
   544 => x"a59b0b80",
   545 => x"f52da590",
   546 => x"0807cc0c",
   547 => x"8ffa0480",
   548 => x"f25182da",
   549 => x"2da59008",
   550 => x"cc0c8fa8",
   551 => x"2da4b008",
   552 => x"982ba590",
   553 => x"08cc0c58",
   554 => x"8fa82da4",
   555 => x"b008902b",
   556 => x"7807a590",
   557 => x"08cc0c58",
   558 => x"8fa82da4",
   559 => x"b008882b",
   560 => x"7807a590",
   561 => x"08cc0c58",
   562 => x"8fa82d77",
   563 => x"a4b00807",
   564 => x"a59008cc",
   565 => x"0c588fa8",
   566 => x"2da4b008",
   567 => x"ff055978",
   568 => x"ff2e80f4",
   569 => x"38a5d457",
   570 => x"79832e80",
   571 => x"f3387652",
   572 => x"77518118",
   573 => x"588de42d",
   574 => x"80ff5676",
   575 => x"70840558",
   576 => x"0870982a",
   577 => x"a5900807",
   578 => x"cc0c558f",
   579 => x"a82d7490",
   580 => x"2a7081ff",
   581 => x"0670a590",
   582 => x"0807cc0c",
   583 => x"51548fa8",
   584 => x"2d74882a",
   585 => x"7081ff06",
   586 => x"70a59008",
   587 => x"07cc0c51",
   588 => x"548fa82d",
   589 => x"7481ff06",
   590 => x"70a59008",
   591 => x"07cc0c55",
   592 => x"8fa82dff",
   593 => x"16567580",
   594 => x"25ffb038",
   595 => x"ff195978",
   596 => x"ff2e0981",
   597 => x"06ff8e38",
   598 => x"a59008cc",
   599 => x"0c8ffa04",
   600 => x"a05182da",
   601 => x"2d775281",
   602 => x"18a9d852",
   603 => x"58a0f92d",
   604 => x"7652a9d8",
   605 => x"51a08b2d",
   606 => x"80ff5691",
   607 => x"fb04a4b0",
   608 => x"0881842e",
   609 => x"bd388184",
   610 => x"0ba4b008",
   611 => x"24fe8038",
   612 => x"a4b00881",
   613 => x"902e8282",
   614 => x"38a4b008",
   615 => x"81fe2e09",
   616 => x"8106fd87",
   617 => x"38a59008",
   618 => x"81fe07cc",
   619 => x"0c8fa82d",
   620 => x"a4b00851",
   621 => x"82da2da5",
   622 => x"900881fe",
   623 => x"07cc0c8f",
   624 => x"fa04a590",
   625 => x"08cc0c8f",
   626 => x"a82da4b0",
   627 => x"08982ba5",
   628 => x"9008cc0c",
   629 => x"588fa82d",
   630 => x"a4b00890",
   631 => x"2b7807a5",
   632 => x"9008cc0c",
   633 => x"588fa82d",
   634 => x"a4b00888",
   635 => x"2b7807a5",
   636 => x"9008cc0c",
   637 => x"588fa82d",
   638 => x"77a4b008",
   639 => x"07a59008",
   640 => x"cc0c588f",
   641 => x"a82da4b0",
   642 => x"085980f7",
   643 => x"5182da2d",
   644 => x"ff195978",
   645 => x"ff2efec0",
   646 => x"38a5d455",
   647 => x"79842e81",
   648 => x"c43880ff",
   649 => x"56a59008",
   650 => x"cc0c8fa8",
   651 => x"2da59008",
   652 => x"cc0ca4b0",
   653 => x"08882b54",
   654 => x"8fa82da5",
   655 => x"9008cc0c",
   656 => x"73a4b008",
   657 => x"07882b54",
   658 => x"8fa82da5",
   659 => x"9008cc0c",
   660 => x"73a4b008",
   661 => x"07882b54",
   662 => x"8fa82d73",
   663 => x"a4b00807",
   664 => x"75708405",
   665 => x"570cff16",
   666 => x"56758025",
   667 => x"ffb73879",
   668 => x"842e8182",
   669 => x"38a5d452",
   670 => x"77518118",
   671 => x"5888872d",
   672 => x"949004a4",
   673 => x"b0088180",
   674 => x"2e098106",
   675 => x"fb9d38a5",
   676 => x"90088180",
   677 => x"07cc0c8f",
   678 => x"fa048056",
   679 => x"a59008cc",
   680 => x"0ca5bc16",
   681 => x"548fa82d",
   682 => x"a4b00874",
   683 => x"81b72d81",
   684 => x"16568b76",
   685 => x"25e63880",
   686 => x"0ba5c70b",
   687 => x"81b72da5",
   688 => x"bc51839e",
   689 => x"2da5bc52",
   690 => x"a9d8519d",
   691 => x"942da4b0",
   692 => x"08802eae",
   693 => x"38a59008",
   694 => x"cc0c8fa8",
   695 => x"2da59008",
   696 => x"cc0c8ffa",
   697 => x"04775281",
   698 => x"18a9d852",
   699 => x"58a0f92d",
   700 => x"80ff5694",
   701 => x"a504a5d4",
   702 => x"52a9d851",
   703 => x"a0c22d94",
   704 => x"9004a590",
   705 => x"0881ff07",
   706 => x"cc0c8fa8",
   707 => x"2da59008",
   708 => x"81ff07cc",
   709 => x"0ca2f051",
   710 => x"839e2d90",
   711 => x"ba0402e8",
   712 => x"050d7779",
   713 => x"7b585555",
   714 => x"80537276",
   715 => x"25a33874",
   716 => x"70810556",
   717 => x"80f52d74",
   718 => x"70810556",
   719 => x"80f52d52",
   720 => x"5271712e",
   721 => x"09810693",
   722 => x"38811353",
   723 => x"757324df",
   724 => x"38800ba4",
   725 => x"b00c0298",
   726 => x"050d0481",
   727 => x"0ba4b00c",
   728 => x"0298050d",
   729 => x"0402d805",
   730 => x"0d800ba9",
   731 => x"fc0ca2f8",
   732 => x"51839e2d",
   733 => x"a5d45280",
   734 => x"518de42d",
   735 => x"a4b00854",
   736 => x"a4b00892",
   737 => x"38a38851",
   738 => x"839e2d73",
   739 => x"5675a4b0",
   740 => x"0c02a805",
   741 => x"0d04a39c",
   742 => x"51839e2d",
   743 => x"8055810b",
   744 => x"a5c80c88",
   745 => x"53a3b452",
   746 => x"a68a5196",
   747 => x"9e2da4b0",
   748 => x"08752e80",
   749 => x"fb388853",
   750 => x"a3c052a6",
   751 => x"a651969e",
   752 => x"2da4b008",
   753 => x"8738a4b0",
   754 => x"08a5c80c",
   755 => x"a5c80880",
   756 => x"2e818938",
   757 => x"a99a0b80",
   758 => x"f52da99b",
   759 => x"0b80f52d",
   760 => x"71982b71",
   761 => x"902b07a9",
   762 => x"9c0b80f5",
   763 => x"2d70882b",
   764 => x"7207a99d",
   765 => x"0b80f52d",
   766 => x"7107a9d2",
   767 => x"0b80f52d",
   768 => x"a9d30b80",
   769 => x"f52d7188",
   770 => x"2b075340",
   771 => x"55525a56",
   772 => x"57557381",
   773 => x"abaa2ea1",
   774 => x"387382d4",
   775 => x"d52ea338",
   776 => x"a3cc5183",
   777 => x"9e2d800b",
   778 => x"a4b00c02",
   779 => x"a8050d04",
   780 => x"a4b008a5",
   781 => x"c80c97b6",
   782 => x"0474518e",
   783 => x"c72da4b0",
   784 => x"0855a5d4",
   785 => x"5274518d",
   786 => x"e42da4b0",
   787 => x"0856a4b0",
   788 => x"08802efe",
   789 => x"b838a3ec",
   790 => x"51839e2d",
   791 => x"8853a3c0",
   792 => x"52a6a651",
   793 => x"969e2da4",
   794 => x"b00881fa",
   795 => x"38810ba9",
   796 => x"fc0ca9d2",
   797 => x"0b80f52d",
   798 => x"547380d5",
   799 => x"2e098106",
   800 => x"ffa438a9",
   801 => x"d30b80f5",
   802 => x"2d547381",
   803 => x"aa2e0981",
   804 => x"06ff9338",
   805 => x"800ba5d4",
   806 => x"0b80f52d",
   807 => x"57547581",
   808 => x"e92e8338",
   809 => x"81547581",
   810 => x"eb2e8c38",
   811 => x"80567376",
   812 => x"2e098106",
   813 => x"fdd738a5",
   814 => x"df0b80f5",
   815 => x"2d5675fe",
   816 => x"e538a5e0",
   817 => x"0b80f52d",
   818 => x"5473822e",
   819 => x"098106fe",
   820 => x"d538a5e1",
   821 => x"0b80f52d",
   822 => x"70aa840c",
   823 => x"ff05a9f8",
   824 => x"0ca5e20b",
   825 => x"80f52da5",
   826 => x"e30b80f5",
   827 => x"2d5b7505",
   828 => x"7a828029",
   829 => x"0570a9ec",
   830 => x"0ca5e40b",
   831 => x"80f52d70",
   832 => x"a9e80ca9",
   833 => x"fc085b59",
   834 => x"577880f8",
   835 => x"38a5e60b",
   836 => x"80f52da5",
   837 => x"e50b80f5",
   838 => x"2d718280",
   839 => x"290570a9",
   840 => x"d40c70a0",
   841 => x"2983ff05",
   842 => x"70892a70",
   843 => x"aa800ca5",
   844 => x"eb0b80f5",
   845 => x"2da5ea0b",
   846 => x"80f52d71",
   847 => x"82802905",
   848 => x"70a5cc0c",
   849 => x"7d71291d",
   850 => x"70a9f40c",
   851 => x"7fa5d00c",
   852 => x"7305aa8c",
   853 => x"0c5a5a51",
   854 => x"51555a81",
   855 => x"5675a4b0",
   856 => x"0c02a805",
   857 => x"0d048853",
   858 => x"a3b452a6",
   859 => x"8a51969e",
   860 => x"2d8056a4",
   861 => x"b008762e",
   862 => x"fdf83875",
   863 => x"a4b00c02",
   864 => x"a8050d04",
   865 => x"8853a3c0",
   866 => x"52a6a651",
   867 => x"969e2da4",
   868 => x"b008fbf9",
   869 => x"38aa8408",
   870 => x"70842ba9",
   871 => x"d40c70aa",
   872 => x"800ca5f9",
   873 => x"0b80f52d",
   874 => x"a5f80b80",
   875 => x"f52d7182",
   876 => x"802905a5",
   877 => x"fa0b80f5",
   878 => x"2d708480",
   879 => x"802912a5",
   880 => x"fb0b80f5",
   881 => x"2d708180",
   882 => x"0a291270",
   883 => x"a5cc0ca9",
   884 => x"e8087129",
   885 => x"a9ec0805",
   886 => x"70aa8c0c",
   887 => x"a6810b80",
   888 => x"f52da680",
   889 => x"0b80f52d",
   890 => x"71828029",
   891 => x"05a6820b",
   892 => x"80f52d70",
   893 => x"84808029",
   894 => x"12a6830b",
   895 => x"80f52d70",
   896 => x"982b81f0",
   897 => x"0a067205",
   898 => x"70a5d00c",
   899 => x"fe117e29",
   900 => x"7705a9f4",
   901 => x"0c525952",
   902 => x"55585e51",
   903 => x"525f525b",
   904 => x"57555781",
   905 => x"569add04",
   906 => x"02ec050d",
   907 => x"7670872c",
   908 => x"7180ff06",
   909 => x"565653a9",
   910 => x"fc088a38",
   911 => x"72882c73",
   912 => x"81ff0655",
   913 => x"55a5d452",
   914 => x"a9ec0815",
   915 => x"518de42d",
   916 => x"a4b00853",
   917 => x"a4b00880",
   918 => x"2e9c38a9",
   919 => x"fc08802e",
   920 => x"9e387310",
   921 => x"10a5d405",
   922 => x"70085253",
   923 => x"8ec72da4",
   924 => x"b008f00a",
   925 => x"065372a4",
   926 => x"b00c0294",
   927 => x"050d0473",
   928 => x"10a5d405",
   929 => x"7080e02d",
   930 => x"52538ef7",
   931 => x"2da4b008",
   932 => x"539cf604",
   933 => x"02cc050d",
   934 => x"7e605d5d",
   935 => x"800ba5d0",
   936 => x"08a9f408",
   937 => x"5a5c57a9",
   938 => x"fc08772e",
   939 => x"818a38aa",
   940 => x"8408842b",
   941 => x"59805675",
   942 => x"792780c4",
   943 => x"38758f06",
   944 => x"a0185854",
   945 => x"73802e80",
   946 => x"fa388077",
   947 => x"80f52d55",
   948 => x"5573752e",
   949 => x"83388155",
   950 => x"7381e52e",
   951 => x"9a388170",
   952 => x"7606555a",
   953 => x"73802e8f",
   954 => x"388b1780",
   955 => x"f52d9806",
   956 => x"5574802e",
   957 => x"80de3881",
   958 => x"16567876",
   959 => x"26ffbe38",
   960 => x"a9fc0880",
   961 => x"2e81c138",
   962 => x"7a519ca8",
   963 => x"2da4b008",
   964 => x"a4b00880",
   965 => x"fffffff8",
   966 => x"06555b73",
   967 => x"80ffffff",
   968 => x"f82e81a4",
   969 => x"38a4b008",
   970 => x"fe05aa84",
   971 => x"0829aa8c",
   972 => x"08055880",
   973 => x"569db704",
   974 => x"aa800884",
   975 => x"2b598056",
   976 => x"9db704a5",
   977 => x"d4527751",
   978 => x"8118588d",
   979 => x"e42da5d4",
   980 => x"579dca04",
   981 => x"8b537b52",
   982 => x"7651969e",
   983 => x"2da4b008",
   984 => x"ff95389c",
   985 => x"1708518e",
   986 => x"c72da4b0",
   987 => x"08841e0c",
   988 => x"9a1780e0",
   989 => x"2d518ef7",
   990 => x"2da4b008",
   991 => x"a4b00855",
   992 => x"56a9fc08",
   993 => x"97387388",
   994 => x"1e0c738c",
   995 => x"1e0c747d",
   996 => x"0c795473",
   997 => x"a4b00c02",
   998 => x"b4050d04",
   999 => x"a4b00888",
  1000 => x"1e0c9417",
  1001 => x"80e02d51",
  1002 => x"8ef72da4",
  1003 => x"b008902b",
  1004 => x"83fff00a",
  1005 => x"06701770",
  1006 => x"7f88050c",
  1007 => x"8c1f0c54",
  1008 => x"747d0c79",
  1009 => x"549f9304",
  1010 => x"800ba4b0",
  1011 => x"0c02b405",
  1012 => x"0d0402f4",
  1013 => x"050d7470",
  1014 => x"08810571",
  1015 => x"0c7008a9",
  1016 => x"f8080653",
  1017 => x"5371802e",
  1018 => x"8b38810b",
  1019 => x"a4b00c02",
  1020 => x"8c050d04",
  1021 => x"88130851",
  1022 => x"9ca82da4",
  1023 => x"b0088814",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba5",
     9 => x"b4080b0b",
    10 => x"0ba5b808",
    11 => x"0b0b0ba5",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a5bc0c0b",
    16 => x"0b0ba5b8",
    17 => x"0c0b0b0b",
    18 => x"a5b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba380",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a5b470ab",
    57 => x"88278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8fd00402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752e80c7",
    65 => x"38875472",
    66 => x"9c2a7384",
    67 => x"2b545271",
    68 => x"802e8338",
    69 => x"81558972",
    70 => x"259938b7",
    71 => x"1252749b",
    72 => x"38ff1454",
    73 => x"738025df",
    74 => x"38800ba5",
    75 => x"b40c0294",
    76 => x"050d04b0",
    77 => x"12527480",
    78 => x"2ee73871",
    79 => x"5182da2d",
    80 => x"ff145473",
    81 => x"8025c038",
    82 => x"82a904b0",
    83 => x"5182da2d",
    84 => x"800ba5b4",
    85 => x"0c029405",
    86 => x"0d0402f8",
    87 => x"050d7352",
    88 => x"c0087088",
    89 => x"2a708106",
    90 => x"51515170",
    91 => x"802ef138",
    92 => x"71c00c71",
    93 => x"a5b40c02",
    94 => x"88050d04",
    95 => x"02f8050d",
    96 => x"7352c408",
    97 => x"70882a70",
    98 => x"81065151",
    99 => x"5170802e",
   100 => x"f13871c4",
   101 => x"0c71a5b4",
   102 => x"0c028805",
   103 => x"0d0402e8",
   104 => x"050d8078",
   105 => x"57557570",
   106 => x"84055708",
   107 => x"53805472",
   108 => x"982a7388",
   109 => x"2b545271",
   110 => x"802ea238",
   111 => x"c0087088",
   112 => x"2a708106",
   113 => x"51515170",
   114 => x"802ef138",
   115 => x"71c00c81",
   116 => x"15811555",
   117 => x"55837425",
   118 => x"d63871ca",
   119 => x"3874a5b4",
   120 => x"0c029805",
   121 => x"0d0402f4",
   122 => x"050dd452",
   123 => x"81ff720c",
   124 => x"71085381",
   125 => x"ff720c72",
   126 => x"882b83fe",
   127 => x"80067208",
   128 => x"7081ff06",
   129 => x"51525381",
   130 => x"ff720c72",
   131 => x"7107882b",
   132 => x"72087081",
   133 => x"ff065152",
   134 => x"5381ff72",
   135 => x"0c727107",
   136 => x"882b7208",
   137 => x"7081ff06",
   138 => x"7207a5b4",
   139 => x"0c525302",
   140 => x"8c050d04",
   141 => x"02f4050d",
   142 => x"74767181",
   143 => x"ff06d40c",
   144 => x"5353a698",
   145 => x"08853871",
   146 => x"892b5271",
   147 => x"982ad40c",
   148 => x"71902a70",
   149 => x"81ff06d4",
   150 => x"0c517188",
   151 => x"2a7081ff",
   152 => x"06d40c51",
   153 => x"7181ff06",
   154 => x"d40c7290",
   155 => x"2a7081ff",
   156 => x"06d40c51",
   157 => x"d4087081",
   158 => x"ff065151",
   159 => x"82b8bf52",
   160 => x"7081ff2e",
   161 => x"09810694",
   162 => x"3881ff0b",
   163 => x"d40cd408",
   164 => x"7081ff06",
   165 => x"ff145451",
   166 => x"5171e538",
   167 => x"70a5b40c",
   168 => x"028c050d",
   169 => x"0402fc05",
   170 => x"0d81c751",
   171 => x"81ff0bd4",
   172 => x"0cff1151",
   173 => x"708025f4",
   174 => x"38028405",
   175 => x"0d0402f0",
   176 => x"050d85a5",
   177 => x"2d819c9f",
   178 => x"53805287",
   179 => x"fc80f751",
   180 => x"84b42da5",
   181 => x"b40854a5",
   182 => x"b408812e",
   183 => x"9038ff13",
   184 => x"5372e638",
   185 => x"72a5b40c",
   186 => x"0290050d",
   187 => x"0481ff0b",
   188 => x"d40c820a",
   189 => x"52849c80",
   190 => x"e95184b4",
   191 => x"2da5b408",
   192 => x"802e8e38",
   193 => x"85a52dff",
   194 => x"135372ff",
   195 => x"bc3885e4",
   196 => x"0481ff0b",
   197 => x"d40c73a5",
   198 => x"b40c0290",
   199 => x"050d0402",
   200 => x"f4050d81",
   201 => x"ff0bd40c",
   202 => x"a3905183",
   203 => x"9e2d9353",
   204 => x"805287fc",
   205 => x"80c15184",
   206 => x"b42da5b4",
   207 => x"08802e93",
   208 => x"3885a52d",
   209 => x"ff135372",
   210 => x"e73872a5",
   211 => x"b40c028c",
   212 => x"050d0481",
   213 => x"ff0bd40c",
   214 => x"810ba5b4",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050d85a5",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"5184b42d",
   221 => x"a5b40881",
   222 => x"2e8f3886",
   223 => x"9f2d8054",
   224 => x"73a5b40c",
   225 => x"0290050d",
   226 => x"0483e62d",
   227 => x"a5b40883",
   228 => x"ffff0653",
   229 => x"7283aa2e",
   230 => x"098106df",
   231 => x"3881ff0b",
   232 => x"d40cb153",
   233 => x"85be2da5",
   234 => x"b4089538",
   235 => x"72822ece",
   236 => x"38ff1353",
   237 => x"72ee3872",
   238 => x"a5b40c02",
   239 => x"90050d04",
   240 => x"805287fc",
   241 => x"80fa5184",
   242 => x"b42da5b4",
   243 => x"08de3881",
   244 => x"ff0bd40c",
   245 => x"d4085381",
   246 => x"ff0bd40c",
   247 => x"81ff0bd4",
   248 => x"0c81ff0b",
   249 => x"d40c81ff",
   250 => x"0bd40c72",
   251 => x"862a7081",
   252 => x"06a5b408",
   253 => x"56515372",
   254 => x"802eff84",
   255 => x"38810ba5",
   256 => x"b40c0290",
   257 => x"050d0402",
   258 => x"e8050d78",
   259 => x"5681ff0b",
   260 => x"d40cd008",
   261 => x"708f2a70",
   262 => x"81065151",
   263 => x"5372f338",
   264 => x"82810bd0",
   265 => x"0c81ff0b",
   266 => x"d40c7752",
   267 => x"87fc80d8",
   268 => x"5184b42d",
   269 => x"a5b40881",
   270 => x"823881ff",
   271 => x"0bd40c81",
   272 => x"fe0bd40c",
   273 => x"80ff5575",
   274 => x"70840557",
   275 => x"0870982a",
   276 => x"d40c7090",
   277 => x"2c7081ff",
   278 => x"06d40c54",
   279 => x"70882c70",
   280 => x"81ff06d4",
   281 => x"0c547081",
   282 => x"ff06d40c",
   283 => x"54ff1555",
   284 => x"748025d3",
   285 => x"3881ff0b",
   286 => x"d40c81ff",
   287 => x"0bd40c81",
   288 => x"ff0bd40c",
   289 => x"868da054",
   290 => x"81ff0bd4",
   291 => x"0cd40881",
   292 => x"ff065574",
   293 => x"8738ff14",
   294 => x"5473ed38",
   295 => x"81ff0bd4",
   296 => x"0cd00870",
   297 => x"8f2a7081",
   298 => x"06515153",
   299 => x"72f33872",
   300 => x"d00c72a5",
   301 => x"b40c0298",
   302 => x"050d04a3",
   303 => x"9451839e",
   304 => x"2d810ba5",
   305 => x"b40c0298",
   306 => x"050d0402",
   307 => x"ec050d76",
   308 => x"78545480",
   309 => x"5580dbc6",
   310 => x"df5281ff",
   311 => x"0bd40cd4",
   312 => x"087081ff",
   313 => x"06515170",
   314 => x"81fe2e95",
   315 => x"38ff1252",
   316 => x"71e83881",
   317 => x"ff0bd40c",
   318 => x"74a5b40c",
   319 => x"0294050d",
   320 => x"04800ba6",
   321 => x"bc0c8373",
   322 => x"259f3883",
   323 => x"e62da5b4",
   324 => x"08747084",
   325 => x"05560ca6",
   326 => x"bc08a5b4",
   327 => x"0805a6bc",
   328 => x"0cfc1353",
   329 => x"728324e3",
   330 => x"38807325",
   331 => x"a03881ff",
   332 => x"0bd40cff",
   333 => x"74708105",
   334 => x"5681b72d",
   335 => x"a6bc0881",
   336 => x"ff05a6bc",
   337 => x"0cff1353",
   338 => x"728024e2",
   339 => x"38815581",
   340 => x"ff0bd40c",
   341 => x"74a5b40c",
   342 => x"0294050d",
   343 => x"0402e805",
   344 => x"0d805287",
   345 => x"fc80c951",
   346 => x"84b42d92",
   347 => x"52a6a851",
   348 => x"89cb2da6",
   349 => x"a80b80f5",
   350 => x"2d81c006",
   351 => x"537280c0",
   352 => x"2e80f738",
   353 => x"a6b10b80",
   354 => x"f52d7010",
   355 => x"8606a6b2",
   356 => x"0b80f52d",
   357 => x"70872a72",
   358 => x"07a6ad0b",
   359 => x"80f52d8f",
   360 => x"06a6ae0b",
   361 => x"80f52d70",
   362 => x"8a2b9880",
   363 => x"06a6af0b",
   364 => x"80f52d70",
   365 => x"822b7207",
   366 => x"a6b00b80",
   367 => x"f52d7086",
   368 => x"2a720782",
   369 => x"1881782b",
   370 => x"81138173",
   371 => x"2b712951",
   372 => x"53585852",
   373 => x"52525259",
   374 => x"53545258",
   375 => x"55558480",
   376 => x"75258e38",
   377 => x"72107581",
   378 => x"2c565374",
   379 => x"848024f4",
   380 => x"3872a5b4",
   381 => x"0c029805",
   382 => x"0d04a6af",
   383 => x"0b80f52d",
   384 => x"a6b00b80",
   385 => x"f52d7190",
   386 => x"2b71882b",
   387 => x"07a6b10b",
   388 => x"80f52d71",
   389 => x"81fffe80",
   390 => x"06077088",
   391 => x"80298880",
   392 => x"05a5b40c",
   393 => x"51555755",
   394 => x"0298050d",
   395 => x"0402f405",
   396 => x"0d810ba6",
   397 => x"980cd008",
   398 => x"708f2a70",
   399 => x"81065151",
   400 => x"5372f338",
   401 => x"72d00c85",
   402 => x"a52da3a4",
   403 => x"51839e2d",
   404 => x"d008708f",
   405 => x"2a708106",
   406 => x"51515372",
   407 => x"f338810b",
   408 => x"d00c8753",
   409 => x"805284d4",
   410 => x"80c05184",
   411 => x"b42da5b4",
   412 => x"08812e8d",
   413 => x"3872822e",
   414 => x"80c538ff",
   415 => x"135372e4",
   416 => x"3886e22d",
   417 => x"a5b408a6",
   418 => x"980ca5b4",
   419 => x"08802eb9",
   420 => x"3881ff0b",
   421 => x"d40c8add",
   422 => x"2da5b408",
   423 => x"a69c0cd0",
   424 => x"08708f2a",
   425 => x"70810651",
   426 => x"515372f3",
   427 => x"3872d00c",
   428 => x"81ff0bd4",
   429 => x"0c810ba5",
   430 => x"b40c028c",
   431 => x"050d0480",
   432 => x"0ba5b40c",
   433 => x"028c050d",
   434 => x"04815287",
   435 => x"fc80d051",
   436 => x"84b42d81",
   437 => x"ff0bd40c",
   438 => x"8add2da5",
   439 => x"b408a69c",
   440 => x"0c8d9f04",
   441 => x"02f0050d",
   442 => x"805481ff",
   443 => x"0bd40cd0",
   444 => x"08708f2a",
   445 => x"70810651",
   446 => x"515372f3",
   447 => x"3882810b",
   448 => x"d00c81ff",
   449 => x"0bd40c75",
   450 => x"5287fc80",
   451 => x"d15184b4",
   452 => x"2da5b408",
   453 => x"802e8a38",
   454 => x"73a5b40c",
   455 => x"0290050d",
   456 => x"04848052",
   457 => x"765189cb",
   458 => x"2da5b408",
   459 => x"54d00870",
   460 => x"8f2a7081",
   461 => x"06515153",
   462 => x"72f33872",
   463 => x"d00c73a5",
   464 => x"b40c0290",
   465 => x"050d0402",
   466 => x"f4050d74",
   467 => x"70882a83",
   468 => x"fe800670",
   469 => x"72982a07",
   470 => x"72882b87",
   471 => x"fc808006",
   472 => x"73982b81",
   473 => x"f00a0671",
   474 => x"730707a5",
   475 => x"b40c5651",
   476 => x"5351028c",
   477 => x"050d0402",
   478 => x"f8050d02",
   479 => x"8e0580f5",
   480 => x"2d74882b",
   481 => x"077083ff",
   482 => x"ff06a5b4",
   483 => x"0c510288",
   484 => x"050d0402",
   485 => x"f8050d73",
   486 => x"70902b71",
   487 => x"902a07a5",
   488 => x"b40c5202",
   489 => x"88050d04",
   490 => x"02f4050d",
   491 => x"a6940853",
   492 => x"cc087082",
   493 => x"80065252",
   494 => x"70732ef4",
   495 => x"38728280",
   496 => x"32a6940c",
   497 => x"71fdff06",
   498 => x"a5b40c02",
   499 => x"8c050d04",
   500 => x"02d8050d",
   501 => x"800ba694",
   502 => x"0ca3a851",
   503 => x"839e2d8c",
   504 => x"ad2d8054",
   505 => x"a5b40874",
   506 => x"2e098106",
   507 => x"8a3873a5",
   508 => x"b40c02a8",
   509 => x"050d04a3",
   510 => x"b051839e",
   511 => x"2d97f02d",
   512 => x"8fa82da5",
   513 => x"b40858a5",
   514 => x"b4088183",
   515 => x"2ebd38a5",
   516 => x"b4088183",
   517 => x"24829238",
   518 => x"a5b40881",
   519 => x"812e82c5",
   520 => x"38a5b408",
   521 => x"81812483",
   522 => x"e138a5b4",
   523 => x"0881802e",
   524 => x"81ec38a3",
   525 => x"b851839e",
   526 => x"2d8fa82d",
   527 => x"a5b40858",
   528 => x"a5b40881",
   529 => x"832e0981",
   530 => x"06c538a6",
   531 => x"9408cc0c",
   532 => x"8fa82da5",
   533 => x"b408982b",
   534 => x"a69408cc",
   535 => x"0c598fa8",
   536 => x"2da5b408",
   537 => x"902b7907",
   538 => x"a69408cc",
   539 => x"0c598fa8",
   540 => x"2da5b408",
   541 => x"882b7907",
   542 => x"a69408cc",
   543 => x"0c598fa8",
   544 => x"2d78a5b4",
   545 => x"0807a694",
   546 => x"08cc0c59",
   547 => x"8fa82da5",
   548 => x"b408ff05",
   549 => x"5a79ff2e",
   550 => x"80fc38a6",
   551 => x"cc577781",
   552 => x"852e85cc",
   553 => x"38765278",
   554 => x"51811959",
   555 => x"8de42d80",
   556 => x"ff567670",
   557 => x"84055808",
   558 => x"55778185",
   559 => x"2e84db38",
   560 => x"74982aa6",
   561 => x"940807cc",
   562 => x"0c8fa82d",
   563 => x"74902a70",
   564 => x"81ff0670",
   565 => x"a6940807",
   566 => x"cc0c5154",
   567 => x"8fa82d74",
   568 => x"882a7081",
   569 => x"ff0670a6",
   570 => x"940807cc",
   571 => x"0c51548f",
   572 => x"a82d7481",
   573 => x"ff0670a6",
   574 => x"940807cc",
   575 => x"0c548fa8",
   576 => x"2dff1656",
   577 => x"758025ff",
   578 => x"a938ff1a",
   579 => x"5a79ff2e",
   580 => x"098106ff",
   581 => x"8638a694",
   582 => x"08cc0c90",
   583 => x"8004a694",
   584 => x"08818007",
   585 => x"cc0c9080",
   586 => x"04a5b408",
   587 => x"81852efe",
   588 => x"9a388185",
   589 => x"0ba5b408",
   590 => x"24829a38",
   591 => x"a5b40881",
   592 => x"fe2e0981",
   593 => x"06fdec38",
   594 => x"a6940881",
   595 => x"fe07cc0c",
   596 => x"8fa82da5",
   597 => x"b4085182",
   598 => x"da2da694",
   599 => x"0881fe07",
   600 => x"cc0c9080",
   601 => x"04a3c051",
   602 => x"839e2da3",
   603 => x"c852aad0",
   604 => x"519e9f2d",
   605 => x"a5b40854",
   606 => x"a5b40880",
   607 => x"2e849b38",
   608 => x"aad40883",
   609 => x"ff05892a",
   610 => x"57805574",
   611 => x"7725fcf0",
   612 => x"38a6cc52",
   613 => x"aad051a1",
   614 => x"962da5b4",
   615 => x"08802e80",
   616 => x"cb38a3d4",
   617 => x"51839e2d",
   618 => x"8056a6cc",
   619 => x"1680f52d",
   620 => x"a6940807",
   621 => x"cc0c8fa8",
   622 => x"2da69408",
   623 => x"802eb838",
   624 => x"ad5182da",
   625 => x"2d811656",
   626 => x"83ff7625",
   627 => x"dd388115",
   628 => x"55747725",
   629 => x"fcaa38aa",
   630 => x"d051a0dd",
   631 => x"2da6cc52",
   632 => x"aad051a1",
   633 => x"962da5b4",
   634 => x"08ffb738",
   635 => x"a5b408a5",
   636 => x"b40c02a8",
   637 => x"050d0480",
   638 => x"df5182da",
   639 => x"2d811656",
   640 => x"83ff7625",
   641 => x"ffa43893",
   642 => x"ce04a3d8",
   643 => x"51839e2d",
   644 => x"a3e052aa",
   645 => x"d0519e9f",
   646 => x"2da69c0b",
   647 => x"80f52da6",
   648 => x"940807cc",
   649 => x"0c8fa82d",
   650 => x"a69d0b80",
   651 => x"f52da694",
   652 => x"0807cc0c",
   653 => x"8fa82da6",
   654 => x"9e0b80f5",
   655 => x"2da69408",
   656 => x"07cc0c8f",
   657 => x"a82da69f",
   658 => x"0b80f52d",
   659 => x"a6940807",
   660 => x"cc0c9080",
   661 => x"04a69408",
   662 => x"cc0c8fa8",
   663 => x"2da5b408",
   664 => x"982ba694",
   665 => x"08cc0c59",
   666 => x"8fa82da5",
   667 => x"b408902b",
   668 => x"7907a694",
   669 => x"08cc0c59",
   670 => x"8fa82da5",
   671 => x"b408882b",
   672 => x"7907a694",
   673 => x"08cc0c59",
   674 => x"8fa82d78",
   675 => x"a5b40807",
   676 => x"a69408cc",
   677 => x"0c598fa8",
   678 => x"2da5b408",
   679 => x"5a905380",
   680 => x"52785181",
   681 => x"f72dff1a",
   682 => x"5a79ff2e",
   683 => x"fce838a6",
   684 => x"cc0ba3ec",
   685 => x"5255839e",
   686 => x"2d80ff56",
   687 => x"a69408cc",
   688 => x"0c8fa82d",
   689 => x"a69408cc",
   690 => x"0ca5b408",
   691 => x"882b548f",
   692 => x"a82da694",
   693 => x"08cc0c73",
   694 => x"a5b40807",
   695 => x"882b548f",
   696 => x"a82da694",
   697 => x"08cc0c73",
   698 => x"a5b40807",
   699 => x"882b548f",
   700 => x"a82d73a5",
   701 => x"b4080775",
   702 => x"70840557",
   703 => x"0cff1656",
   704 => x"758025ff",
   705 => x"b738a3ec",
   706 => x"51839e2d",
   707 => x"a6cc5278",
   708 => x"51811959",
   709 => x"88872d95",
   710 => x"a6049053",
   711 => x"80527451",
   712 => x"81f72d74",
   713 => x"982aa694",
   714 => x"0807cc0c",
   715 => x"8fa82d74",
   716 => x"902a7081",
   717 => x"ff0670a6",
   718 => x"940807cc",
   719 => x"0c51548f",
   720 => x"a82d7488",
   721 => x"2a7081ff",
   722 => x"0670a694",
   723 => x"0807cc0c",
   724 => x"51548fa8",
   725 => x"2d7481ff",
   726 => x"0670a694",
   727 => x"0807cc0c",
   728 => x"548fa82d",
   729 => x"ff165675",
   730 => x"8025fac6",
   731 => x"38928a04",
   732 => x"a3f05183",
   733 => x"9e2d9053",
   734 => x"80527851",
   735 => x"81f72da0",
   736 => x"5182da2d",
   737 => x"7852aad0",
   738 => x"51a1cd2d",
   739 => x"7652aad0",
   740 => x"51a1962d",
   741 => x"80ff5691",
   742 => x"b204a3f4",
   743 => x"51839e2d",
   744 => x"73a5b40c",
   745 => x"02a8050d",
   746 => x"0402e805",
   747 => x"0d77797b",
   748 => x"58555580",
   749 => x"53727625",
   750 => x"a3387470",
   751 => x"81055680",
   752 => x"f52d7470",
   753 => x"81055680",
   754 => x"f52d5252",
   755 => x"71712e09",
   756 => x"81069338",
   757 => x"81135375",
   758 => x"7324df38",
   759 => x"800ba5b4",
   760 => x"0c029805",
   761 => x"0d04810b",
   762 => x"a5b40c02",
   763 => x"98050d04",
   764 => x"02d8050d",
   765 => x"800baaf4",
   766 => x"0ca3fc51",
   767 => x"839e2da6",
   768 => x"cc528051",
   769 => x"8de42da5",
   770 => x"b40854a5",
   771 => x"b4089238",
   772 => x"a48c5183",
   773 => x"9e2d7356",
   774 => x"75a5b40c",
   775 => x"02a8050d",
   776 => x"04a4a051",
   777 => x"839e2d80",
   778 => x"55810ba6",
   779 => x"c00c8853",
   780 => x"a4b852a7",
   781 => x"825197a9",
   782 => x"2da5b408",
   783 => x"752e80fb",
   784 => x"388853a4",
   785 => x"c452a79e",
   786 => x"5197a92d",
   787 => x"a5b40887",
   788 => x"38a5b408",
   789 => x"a6c00ca6",
   790 => x"c008802e",
   791 => x"818938aa",
   792 => x"920b80f5",
   793 => x"2daa930b",
   794 => x"80f52d71",
   795 => x"982b7190",
   796 => x"2b07aa94",
   797 => x"0b80f52d",
   798 => x"70882b72",
   799 => x"07aa950b",
   800 => x"80f52d71",
   801 => x"07aaca0b",
   802 => x"80f52daa",
   803 => x"cb0b80f5",
   804 => x"2d71882b",
   805 => x"07534055",
   806 => x"525a5657",
   807 => x"557381ab",
   808 => x"aa2ea138",
   809 => x"7382d4d5",
   810 => x"2ea338a4",
   811 => x"d051839e",
   812 => x"2d800ba5",
   813 => x"b40c02a8",
   814 => x"050d04a5",
   815 => x"b408a6c0",
   816 => x"0c98c104",
   817 => x"74518ec7",
   818 => x"2da5b408",
   819 => x"55a6cc52",
   820 => x"74518de4",
   821 => x"2da5b408",
   822 => x"56a5b408",
   823 => x"802efeb8",
   824 => x"38a4f051",
   825 => x"839e2d88",
   826 => x"53a4c452",
   827 => x"a79e5197",
   828 => x"a92da5b4",
   829 => x"0881fa38",
   830 => x"810baaf4",
   831 => x"0caaca0b",
   832 => x"80f52d54",
   833 => x"7380d52e",
   834 => x"098106ff",
   835 => x"a438aacb",
   836 => x"0b80f52d",
   837 => x"547381aa",
   838 => x"2e098106",
   839 => x"ff933880",
   840 => x"0ba6cc0b",
   841 => x"80f52d57",
   842 => x"547581e9",
   843 => x"2e833881",
   844 => x"547581eb",
   845 => x"2e8c3880",
   846 => x"5673762e",
   847 => x"098106fd",
   848 => x"d738a6d7",
   849 => x"0b80f52d",
   850 => x"5675fee5",
   851 => x"38a6d80b",
   852 => x"80f52d54",
   853 => x"73822e09",
   854 => x"8106fed5",
   855 => x"38a6d90b",
   856 => x"80f52d70",
   857 => x"aafc0cff",
   858 => x"05aaf00c",
   859 => x"a6da0b80",
   860 => x"f52da6db",
   861 => x"0b80f52d",
   862 => x"5b75057a",
   863 => x"82802905",
   864 => x"70aae40c",
   865 => x"a6dc0b80",
   866 => x"f52d70aa",
   867 => x"e00caaf4",
   868 => x"085b5957",
   869 => x"7880f838",
   870 => x"a6de0b80",
   871 => x"f52da6dd",
   872 => x"0b80f52d",
   873 => x"71828029",
   874 => x"0570aacc",
   875 => x"0c70a029",
   876 => x"83ff0570",
   877 => x"892a70aa",
   878 => x"f80ca6e3",
   879 => x"0b80f52d",
   880 => x"a6e20b80",
   881 => x"f52d7182",
   882 => x"80290570",
   883 => x"a6c40c7d",
   884 => x"71291d70",
   885 => x"aaec0c7f",
   886 => x"a6c80c73",
   887 => x"05ab840c",
   888 => x"5a5a5151",
   889 => x"555a8156",
   890 => x"75a5b40c",
   891 => x"02a8050d",
   892 => x"048853a4",
   893 => x"b852a782",
   894 => x"5197a92d",
   895 => x"8056a5b4",
   896 => x"08762efd",
   897 => x"f83875a5",
   898 => x"b40c02a8",
   899 => x"050d0488",
   900 => x"53a4c452",
   901 => x"a79e5197",
   902 => x"a92da5b4",
   903 => x"08fbf938",
   904 => x"aafc0870",
   905 => x"842baacc",
   906 => x"0c70aaf8",
   907 => x"0ca6f10b",
   908 => x"80f52da6",
   909 => x"f00b80f5",
   910 => x"2d718280",
   911 => x"2905a6f2",
   912 => x"0b80f52d",
   913 => x"70848080",
   914 => x"2912a6f3",
   915 => x"0b80f52d",
   916 => x"7081800a",
   917 => x"291270a6",
   918 => x"c40caae0",
   919 => x"087129aa",
   920 => x"e4080570",
   921 => x"ab840ca6",
   922 => x"f90b80f5",
   923 => x"2da6f80b",
   924 => x"80f52d71",
   925 => x"82802905",
   926 => x"a6fa0b80",
   927 => x"f52d7084",
   928 => x"80802912",
   929 => x"a6fb0b80",
   930 => x"f52d7098",
   931 => x"2b81f00a",
   932 => x"06720570",
   933 => x"a6c80cfe",
   934 => x"117e2977",
   935 => x"05aaec0c",
   936 => x"52595255",
   937 => x"585e5152",
   938 => x"5f525b57",
   939 => x"55578156",
   940 => x"9be80402",
   941 => x"ec050d76",
   942 => x"70872c71",
   943 => x"80ff0656",
   944 => x"5653aaf4",
   945 => x"088a3872",
   946 => x"882c7381",
   947 => x"ff065555",
   948 => x"a6cc52aa",
   949 => x"e4081551",
   950 => x"8de42da5",
   951 => x"b40853a5",
   952 => x"b408802e",
   953 => x"9c38aaf4",
   954 => x"08802e9e",
   955 => x"38731010",
   956 => x"a6cc0570",
   957 => x"0852538e",
   958 => x"c72da5b4",
   959 => x"08f00a06",
   960 => x"5372a5b4",
   961 => x"0c029405",
   962 => x"0d047310",
   963 => x"a6cc0570",
   964 => x"80e02d52",
   965 => x"538ef72d",
   966 => x"a5b40853",
   967 => x"9e810402",
   968 => x"cc050d7e",
   969 => x"605d5d80",
   970 => x"0ba6c808",
   971 => x"aaec085a",
   972 => x"5c57aaf4",
   973 => x"08772e81",
   974 => x"8a38aafc",
   975 => x"08842b59",
   976 => x"80567579",
   977 => x"2780c438",
   978 => x"758f06a0",
   979 => x"18585473",
   980 => x"802e80fa",
   981 => x"38807780",
   982 => x"f52d5555",
   983 => x"73752e83",
   984 => x"38815573",
   985 => x"81e52e9a",
   986 => x"38817076",
   987 => x"06555a73",
   988 => x"802e8f38",
   989 => x"8b1780f5",
   990 => x"2d980655",
   991 => x"74802e80",
   992 => x"de388116",
   993 => x"56787626",
   994 => x"ffbe38aa",
   995 => x"f408802e",
   996 => x"81c1387a",
   997 => x"519db32d",
   998 => x"a5b408a5",
   999 => x"b40880ff",
  1000 => x"fffff806",
  1001 => x"555b7380",
  1002 => x"fffffff8",
  1003 => x"2e81a438",
  1004 => x"a5b408fe",
  1005 => x"05aafc08",
  1006 => x"29ab8408",
  1007 => x"05588056",
  1008 => x"9ec204aa",
  1009 => x"f808842b",
  1010 => x"5980569e",
  1011 => x"c204a6cc",
  1012 => x"52775181",
  1013 => x"18588de4",
  1014 => x"2da6cc57",
  1015 => x"9ed5048b",
  1016 => x"537b5276",
  1017 => x"5197a92d",
  1018 => x"a5b408ff",
  1019 => x"95389c17",
  1020 => x"08518ec7",
  1021 => x"2da5b408",
  1022 => x"841e0c9a",
  1023 => x"1780e02d",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0b9e",
     9 => x"f8080b0b",
    10 => x"0b9efc08",
    11 => x"0b0b0b9f",
    12 => x"80080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"9f800c0b",
    16 => x"0b0b9efc",
    17 => x"0c0b0b0b",
    18 => x"9ef80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b9bb0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"9ef870a3",
    57 => x"f8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"90b10402",
    62 => x"f8050d73",
    63 => x"52c00870",
    64 => x"882a7081",
    65 => x"06515151",
    66 => x"70802ef1",
    67 => x"3871c00c",
    68 => x"719ef80c",
    69 => x"0288050d",
    70 => x"0402f805",
    71 => x"0d7352c4",
    72 => x"0870882a",
    73 => x"70810651",
    74 => x"51517080",
    75 => x"2ef13871",
    76 => x"c40c719e",
    77 => x"f80c0288",
    78 => x"050d0402",
    79 => x"e8050d80",
    80 => x"78575575",
    81 => x"70840557",
    82 => x"08538054",
    83 => x"72982a73",
    84 => x"882b5452",
    85 => x"71802ea2",
    86 => x"38c00870",
    87 => x"882a7081",
    88 => x"06515151",
    89 => x"70802ef1",
    90 => x"3871c00c",
    91 => x"81158115",
    92 => x"55558374",
    93 => x"25d63871",
    94 => x"ca38749e",
    95 => x"f80c0298",
    96 => x"050d0402",
    97 => x"f4050dd4",
    98 => x"5281ff72",
    99 => x"0c710853",
   100 => x"81ff720c",
   101 => x"72882b83",
   102 => x"fe800672",
   103 => x"087081ff",
   104 => x"06515253",
   105 => x"81ff720c",
   106 => x"72710788",
   107 => x"2b720870",
   108 => x"81ff0651",
   109 => x"525381ff",
   110 => x"720c7271",
   111 => x"07882b72",
   112 => x"087081ff",
   113 => x"0672079e",
   114 => x"f80c5253",
   115 => x"028c050d",
   116 => x"0402f405",
   117 => x"0d747671",
   118 => x"81ff06d4",
   119 => x"0c53539f",
   120 => x"8c088538",
   121 => x"71892b52",
   122 => x"71982ad4",
   123 => x"0c71902a",
   124 => x"7081ff06",
   125 => x"d40c5171",
   126 => x"882a7081",
   127 => x"ff06d40c",
   128 => x"517181ff",
   129 => x"06d40c72",
   130 => x"902a7081",
   131 => x"ff06d40c",
   132 => x"51d40870",
   133 => x"81ff0651",
   134 => x"5182b8bf",
   135 => x"527081ff",
   136 => x"2e098106",
   137 => x"943881ff",
   138 => x"0bd40cd4",
   139 => x"087081ff",
   140 => x"06ff1454",
   141 => x"515171e5",
   142 => x"38709ef8",
   143 => x"0c028c05",
   144 => x"0d0402fc",
   145 => x"050d81c7",
   146 => x"5181ff0b",
   147 => x"d40cff11",
   148 => x"51708025",
   149 => x"f4380284",
   150 => x"050d0402",
   151 => x"f0050d84",
   152 => x"c22d819c",
   153 => x"9f538052",
   154 => x"87fc80f7",
   155 => x"5183d12d",
   156 => x"9ef80854",
   157 => x"9ef80881",
   158 => x"2e098106",
   159 => x"a33881ff",
   160 => x"0bd40c82",
   161 => x"0a52849c",
   162 => x"80e95183",
   163 => x"d12d9ef8",
   164 => x"088b3881",
   165 => x"ff0bd40c",
   166 => x"735385a6",
   167 => x"0484c22d",
   168 => x"ff135372",
   169 => x"c138729e",
   170 => x"f80c0290",
   171 => x"050d0402",
   172 => x"f4050d81",
   173 => x"ff0bd40c",
   174 => x"9bc05182",
   175 => x"bb2d9353",
   176 => x"805287fc",
   177 => x"80c15183",
   178 => x"d12d9ef8",
   179 => x"088b3881",
   180 => x"ff0bd40c",
   181 => x"815385e2",
   182 => x"0484c22d",
   183 => x"ff135372",
   184 => x"df38729e",
   185 => x"f80c028c",
   186 => x"050d0402",
   187 => x"f0050d84",
   188 => x"c22d83aa",
   189 => x"52849c80",
   190 => x"c85183d1",
   191 => x"2d9ef808",
   192 => x"812e0981",
   193 => x"06923883",
   194 => x"832d9ef8",
   195 => x"0883ffff",
   196 => x"06537283",
   197 => x"aa2e9138",
   198 => x"85af2d86",
   199 => x"a3048154",
   200 => x"87880480",
   201 => x"54878804",
   202 => x"81ff0bd4",
   203 => x"0cb15384",
   204 => x"db2d9ef8",
   205 => x"08802e80",
   206 => x"c0388052",
   207 => x"87fc80fa",
   208 => x"5183d12d",
   209 => x"9ef808b1",
   210 => x"3881ff0b",
   211 => x"d40cd408",
   212 => x"5381ff0b",
   213 => x"d40c81ff",
   214 => x"0bd40c81",
   215 => x"ff0bd40c",
   216 => x"81ff0bd4",
   217 => x"0c72862a",
   218 => x"7081069e",
   219 => x"f8085651",
   220 => x"5372802e",
   221 => x"9338869e",
   222 => x"0472822e",
   223 => x"ffa538ff",
   224 => x"135372ff",
   225 => x"aa387254",
   226 => x"739ef80c",
   227 => x"0290050d",
   228 => x"04800b9e",
   229 => x"f80c0402",
   230 => x"ec050d76",
   231 => x"78535480",
   232 => x"5580dbc6",
   233 => x"df5381ff",
   234 => x"0bd40cd4",
   235 => x"087081ff",
   236 => x"06515170",
   237 => x"81fe2e09",
   238 => x"810680ce",
   239 => x"38800b9f",
   240 => x"b00c8372",
   241 => x"259d3883",
   242 => x"832d9ef8",
   243 => x"08747084",
   244 => x"05560c9f",
   245 => x"b0089ef8",
   246 => x"08059fb0",
   247 => x"0cfc1252",
   248 => x"87c20480",
   249 => x"72259e38",
   250 => x"81ff0bd4",
   251 => x"0cff7470",
   252 => x"81055681",
   253 => x"b72d9fb0",
   254 => x"0881ff05",
   255 => x"9fb00cff",
   256 => x"125287e3",
   257 => x"04815588",
   258 => x"9104ff13",
   259 => x"5372ff96",
   260 => x"3881ff0b",
   261 => x"d40c749e",
   262 => x"f80c0294",
   263 => x"050d0402",
   264 => x"e8050d80",
   265 => x"5287fc80",
   266 => x"c95183d1",
   267 => x"2d92529f",
   268 => x"9c518797",
   269 => x"2d9f9c0b",
   270 => x"80f52d81",
   271 => x"c0065372",
   272 => x"80c02e09",
   273 => x"8106b038",
   274 => x"9fa30b80",
   275 => x"f52d9fa4",
   276 => x"0b80f52d",
   277 => x"71902b71",
   278 => x"882b079f",
   279 => x"a50b80f5",
   280 => x"2d7181ff",
   281 => x"fe800607",
   282 => x"70888029",
   283 => x"88800551",
   284 => x"51555755",
   285 => x"89e1049f",
   286 => x"a50b80f5",
   287 => x"2d701086",
   288 => x"069fa60b",
   289 => x"80f52d70",
   290 => x"872a7207",
   291 => x"9fa10b80",
   292 => x"f52d8f06",
   293 => x"9fa20b80",
   294 => x"f52d708a",
   295 => x"2b988006",
   296 => x"9fa30b80",
   297 => x"f52d7082",
   298 => x"2b72079f",
   299 => x"a40b80f5",
   300 => x"2d70862a",
   301 => x"72078218",
   302 => x"81782b81",
   303 => x"1381732b",
   304 => x"71295153",
   305 => x"58585252",
   306 => x"52525953",
   307 => x"54525855",
   308 => x"55848075",
   309 => x"258b3872",
   310 => x"1075812c",
   311 => x"565389d1",
   312 => x"04729ef8",
   313 => x"0c029805",
   314 => x"0d0402f4",
   315 => x"050d810b",
   316 => x"9f8c0cd0",
   317 => x"08708f2a",
   318 => x"70810651",
   319 => x"515372f3",
   320 => x"3872d00c",
   321 => x"84c22d9b",
   322 => x"c45182bb",
   323 => x"2dd00870",
   324 => x"8f2a7081",
   325 => x"06515153",
   326 => x"72f33881",
   327 => x"0bd00c87",
   328 => x"53805284",
   329 => x"d480c051",
   330 => x"83d12d9e",
   331 => x"f808812e",
   332 => x"94387282",
   333 => x"2e098106",
   334 => x"86388053",
   335 => x"8b8304ff",
   336 => x"135372dd",
   337 => x"3885eb2d",
   338 => x"9ef8089f",
   339 => x"8c0c9ef8",
   340 => x"088b3881",
   341 => x"5287fc80",
   342 => x"d05183d1",
   343 => x"2d81ff0b",
   344 => x"d40c889f",
   345 => x"2d9ef808",
   346 => x"9f900cd0",
   347 => x"08708f2a",
   348 => x"70810651",
   349 => x"515372f3",
   350 => x"3872d00c",
   351 => x"81ff0bd4",
   352 => x"0c815372",
   353 => x"9ef80c02",
   354 => x"8c050d04",
   355 => x"02f0050d",
   356 => x"805481ff",
   357 => x"0bd40cd0",
   358 => x"08708f2a",
   359 => x"70810651",
   360 => x"515372f3",
   361 => x"3882810b",
   362 => x"d00c81ff",
   363 => x"0bd40c75",
   364 => x"5287fc80",
   365 => x"d15183d1",
   366 => x"2d9ef808",
   367 => x"9e388480",
   368 => x"52765187",
   369 => x"972d9ef8",
   370 => x"0854d008",
   371 => x"708f2a70",
   372 => x"81065151",
   373 => x"5372f338",
   374 => x"72d00c73",
   375 => x"9ef80c02",
   376 => x"90050d04",
   377 => x"02f4050d",
   378 => x"7470882a",
   379 => x"83fe8006",
   380 => x"7072982a",
   381 => x"0772882b",
   382 => x"87fc8080",
   383 => x"0673982b",
   384 => x"81f00a06",
   385 => x"71730707",
   386 => x"9ef80c56",
   387 => x"51535102",
   388 => x"8c050d04",
   389 => x"02f8050d",
   390 => x"028e0580",
   391 => x"f52d7488",
   392 => x"2b077083",
   393 => x"ffff069e",
   394 => x"f80c5102",
   395 => x"88050d04",
   396 => x"02f8050d",
   397 => x"7370902b",
   398 => x"71902a07",
   399 => x"9ef80c52",
   400 => x"0288050d",
   401 => x"0402f405",
   402 => x"0d9f8808",
   403 => x"53cc0870",
   404 => x"82800652",
   405 => x"5270732e",
   406 => x"f4387282",
   407 => x"80329f88",
   408 => x"0c71fdff",
   409 => x"069ef80c",
   410 => x"028c050d",
   411 => x"0402e005",
   412 => x"0d795780",
   413 => x"0b9f880c",
   414 => x"8cc52d9e",
   415 => x"f808539e",
   416 => x"f8088181",
   417 => x"2e828d38",
   418 => x"9ef80881",
   419 => x"81248c38",
   420 => x"9ef80881",
   421 => x"802e9838",
   422 => x"9098049e",
   423 => x"f8088182",
   424 => x"2e81ad38",
   425 => x"9ef80881",
   426 => x"832e9338",
   427 => x"9098049b",
   428 => x"cc5182bb",
   429 => x"2d9f8808",
   430 => x"7307538f",
   431 => x"8e049bc8",
   432 => x"5182bb2d",
   433 => x"9f8808cc",
   434 => x"0c8cc52d",
   435 => x"9ef80898",
   436 => x"2b9f8808",
   437 => x"cc0c548c",
   438 => x"c52d9ef8",
   439 => x"08902b74",
   440 => x"079f8808",
   441 => x"cc0c548c",
   442 => x"c52d9ef8",
   443 => x"08882b74",
   444 => x"079f8808",
   445 => x"cc0c548c",
   446 => x"c52d739e",
   447 => x"f808079f",
   448 => x"8808cc0c",
   449 => x"548cc52d",
   450 => x"9ef8089b",
   451 => x"d8525682",
   452 => x"bb2dff16",
   453 => x"5675ff2e",
   454 => x"af389fc0",
   455 => x"52735181",
   456 => x"14548b8c",
   457 => x"2d9bec51",
   458 => x"82bb2d80",
   459 => x"559fc015",
   460 => x"80f52d9f",
   461 => x"880807cc",
   462 => x"0c8cc52d",
   463 => x"81155583",
   464 => x"ff7525e9",
   465 => x"388e9204",
   466 => x"9f8808cc",
   467 => x"0c909e04",
   468 => x"9bfc5182",
   469 => x"bb2d9f90",
   470 => x"0b80f52d",
   471 => x"9f880807",
   472 => x"cc0c8cc5",
   473 => x"2d9f910b",
   474 => x"80f52d9f",
   475 => x"880807cc",
   476 => x"0c8cc52d",
   477 => x"9f920b80",
   478 => x"f52d9f88",
   479 => x"0807cc0c",
   480 => x"8cc52d9f",
   481 => x"930b80f5",
   482 => x"2d9f8808",
   483 => x"075372cc",
   484 => x"0c909e04",
   485 => x"9c905182",
   486 => x"bb2d7652",
   487 => x"a3c45197",
   488 => x"d32d9ef8",
   489 => x"08802e80",
   490 => x"e638a3c8",
   491 => x"0883ff05",
   492 => x"892a5680",
   493 => x"54737625",
   494 => x"80e4389f",
   495 => x"c052a3c4",
   496 => x"519a982d",
   497 => x"9ef80880",
   498 => x"2e80dc38",
   499 => x"9bec5182",
   500 => x"bb2d8055",
   501 => x"9fc01580",
   502 => x"f52d9f88",
   503 => x"0807cc0c",
   504 => x"8cc52d9f",
   505 => x"8808802e",
   506 => x"8638ad51",
   507 => x"8ff20480",
   508 => x"df5181f7",
   509 => x"2d811555",
   510 => x"83ff7525",
   511 => x"d7388114",
   512 => x"54737625",
   513 => x"9938a3c4",
   514 => x"5199eb2d",
   515 => x"8fbb049c",
   516 => x"a05182bb",
   517 => x"2d90a704",
   518 => x"9cb45182",
   519 => x"bb2d9cc8",
   520 => x"5182bb2d",
   521 => x"8cf80480",
   522 => x"0b9ef80c",
   523 => x"02a0050d",
   524 => x"0402fc05",
   525 => x"0d9ce451",
   526 => x"82bb2d89",
   527 => x"ea2d9ef8",
   528 => x"08802ea3",
   529 => x"389cfc51",
   530 => x"82bb2d91",
   531 => x"af2d9d94",
   532 => x"518ced2d",
   533 => x"9ef80880",
   534 => x"2e87389d",
   535 => x"a05190e4",
   536 => x"049dac51",
   537 => x"82bb2d80",
   538 => x"0b9ef80c",
   539 => x"0284050d",
   540 => x"0402e805",
   541 => x"0d77797b",
   542 => x"58555580",
   543 => x"53727625",
   544 => x"a3387470",
   545 => x"81055680",
   546 => x"f52d7470",
   547 => x"81055680",
   548 => x"f52d5252",
   549 => x"71712e86",
   550 => x"38815191",
   551 => x"a6048113",
   552 => x"5390fd04",
   553 => x"8051709e",
   554 => x"f80c0298",
   555 => x"050d0402",
   556 => x"d8050d80",
   557 => x"0ba3e40c",
   558 => x"9dc05182",
   559 => x"bb2d9fc0",
   560 => x"5280518b",
   561 => x"8c2d9ef8",
   562 => x"08549ef8",
   563 => x"088c389d",
   564 => x"d05182bb",
   565 => x"2d735596",
   566 => x"dc049de4",
   567 => x"5182bb2d",
   568 => x"8056810b",
   569 => x"9fb40c88",
   570 => x"539dfc52",
   571 => x"9ff65190",
   572 => x"f12d9ef8",
   573 => x"08762e09",
   574 => x"81068738",
   575 => x"9ef8089f",
   576 => x"b40c8853",
   577 => x"9e8852a0",
   578 => x"925190f1",
   579 => x"2d9ef808",
   580 => x"87389ef8",
   581 => x"089fb40c",
   582 => x"9fb40880",
   583 => x"2e80ff38",
   584 => x"a3860b80",
   585 => x"f52da387",
   586 => x"0b80f52d",
   587 => x"71982b71",
   588 => x"902b07a3",
   589 => x"880b80f5",
   590 => x"2d70882b",
   591 => x"7207a389",
   592 => x"0b80f52d",
   593 => x"7107a3be",
   594 => x"0b80f52d",
   595 => x"a3bf0b80",
   596 => x"f52d7188",
   597 => x"2b07535f",
   598 => x"54525a56",
   599 => x"57557381",
   600 => x"abaa2e09",
   601 => x"81068d38",
   602 => x"75518be4",
   603 => x"2d9ef808",
   604 => x"56938404",
   605 => x"7382d4d5",
   606 => x"2e8a389e",
   607 => x"945182bb",
   608 => x"2d94a804",
   609 => x"9fc05275",
   610 => x"518b8c2d",
   611 => x"9ef80855",
   612 => x"9ef80880",
   613 => x"2e83c538",
   614 => x"9eb45182",
   615 => x"bb2d8853",
   616 => x"9e8852a0",
   617 => x"925190f1",
   618 => x"2d9ef808",
   619 => x"8938810b",
   620 => x"a3e40c93",
   621 => x"ce048853",
   622 => x"9dfc529f",
   623 => x"f65190f1",
   624 => x"2d80559e",
   625 => x"f808752e",
   626 => x"09810683",
   627 => x"8f38a3be",
   628 => x"0b80f52d",
   629 => x"547380d5",
   630 => x"2e098106",
   631 => x"80ca38a3",
   632 => x"bf0b80f5",
   633 => x"2d547381",
   634 => x"aa2e0981",
   635 => x"06ba3880",
   636 => x"0b9fc00b",
   637 => x"80f52d56",
   638 => x"547481e9",
   639 => x"2e833881",
   640 => x"547481eb",
   641 => x"2e8c3880",
   642 => x"5573752e",
   643 => x"09810682",
   644 => x"cb389fcb",
   645 => x"0b80f52d",
   646 => x"55748d38",
   647 => x"9fcc0b80",
   648 => x"f52d5473",
   649 => x"822e8638",
   650 => x"805596dc",
   651 => x"049fcd0b",
   652 => x"80f52d70",
   653 => x"a3ec0cff",
   654 => x"05a3e00c",
   655 => x"9fce0b80",
   656 => x"f52d9fcf",
   657 => x"0b80f52d",
   658 => x"58760577",
   659 => x"82802905",
   660 => x"70a3d40c",
   661 => x"9fd00b80",
   662 => x"f52d70a3",
   663 => x"d00ca3e4",
   664 => x"08595758",
   665 => x"76802e81",
   666 => x"a3388853",
   667 => x"9e8852a0",
   668 => x"925190f1",
   669 => x"2d9ef808",
   670 => x"81e238a3",
   671 => x"ec087084",
   672 => x"2ba3c00c",
   673 => x"70a3e80c",
   674 => x"9fe50b80",
   675 => x"f52d9fe4",
   676 => x"0b80f52d",
   677 => x"71828029",
   678 => x"059fe60b",
   679 => x"80f52d70",
   680 => x"84808029",
   681 => x"129fe70b",
   682 => x"80f52d70",
   683 => x"81800a29",
   684 => x"12709fb8",
   685 => x"0ca3d008",
   686 => x"7129a3d4",
   687 => x"080570a3",
   688 => x"f40c9fed",
   689 => x"0b80f52d",
   690 => x"9fec0b80",
   691 => x"f52d7182",
   692 => x"8029059f",
   693 => x"ee0b80f5",
   694 => x"2d708480",
   695 => x"8029129f",
   696 => x"ef0b80f5",
   697 => x"2d70982b",
   698 => x"81f00a06",
   699 => x"7205709f",
   700 => x"bc0cfe11",
   701 => x"7e297705",
   702 => x"a3dc0c52",
   703 => x"59524354",
   704 => x"5e515259",
   705 => x"525d5759",
   706 => x"5796da04",
   707 => x"9fd20b80",
   708 => x"f52d9fd1",
   709 => x"0b80f52d",
   710 => x"71828029",
   711 => x"0570a3c0",
   712 => x"0c70a029",
   713 => x"83ff0570",
   714 => x"892a70a3",
   715 => x"e80c9fd7",
   716 => x"0b80f52d",
   717 => x"9fd60b80",
   718 => x"f52d7182",
   719 => x"80290570",
   720 => x"9fb80c7b",
   721 => x"71291e70",
   722 => x"a3dc0c7d",
   723 => x"9fbc0c73",
   724 => x"05a3f40c",
   725 => x"555e5151",
   726 => x"55558155",
   727 => x"749ef80c",
   728 => x"02a8050d",
   729 => x"0402ec05",
   730 => x"0d767087",
   731 => x"2c7180ff",
   732 => x"06555654",
   733 => x"a3e4088a",
   734 => x"3873882c",
   735 => x"7481ff06",
   736 => x"54559fc0",
   737 => x"52a3d408",
   738 => x"15518b8c",
   739 => x"2d9ef808",
   740 => x"549ef808",
   741 => x"802eb338",
   742 => x"a3e40880",
   743 => x"2e983872",
   744 => x"84299fc0",
   745 => x"05700852",
   746 => x"538be42d",
   747 => x"9ef808f0",
   748 => x"0a065397",
   749 => x"c8047210",
   750 => x"9fc00570",
   751 => x"80e02d52",
   752 => x"538c942d",
   753 => x"9ef80853",
   754 => x"7254739e",
   755 => x"f80c0294",
   756 => x"050d0402",
   757 => x"c8050d7f",
   758 => x"615f5b80",
   759 => x"0b9fbc08",
   760 => x"a3dc0859",
   761 => x"5d56a3e4",
   762 => x"08762e8a",
   763 => x"38a3ec08",
   764 => x"842b5897",
   765 => x"fc04a3e8",
   766 => x"08842b58",
   767 => x"80597878",
   768 => x"2781a938",
   769 => x"788f06a0",
   770 => x"17575473",
   771 => x"8f389fc0",
   772 => x"52765181",
   773 => x"17578b8c",
   774 => x"2d9fc056",
   775 => x"807680f5",
   776 => x"2d565474",
   777 => x"742e8338",
   778 => x"81547481",
   779 => x"e52e80f6",
   780 => x"38817075",
   781 => x"06555d73",
   782 => x"802e80ea",
   783 => x"388b1680",
   784 => x"f52d9806",
   785 => x"5a7980de",
   786 => x"388b537d",
   787 => x"52755190",
   788 => x"f12d9ef8",
   789 => x"0880cf38",
   790 => x"9c160851",
   791 => x"8be42d9e",
   792 => x"f808841c",
   793 => x"0c9a1680",
   794 => x"e02d518c",
   795 => x"942d9ef8",
   796 => x"089ef808",
   797 => x"881d0c9e",
   798 => x"f8085555",
   799 => x"a3e40880",
   800 => x"2e983894",
   801 => x"1680e02d",
   802 => x"518c942d",
   803 => x"9ef80890",
   804 => x"2b83fff0",
   805 => x"0a067016",
   806 => x"51547388",
   807 => x"1c0c797b",
   808 => x"0c7c5499",
   809 => x"e2048119",
   810 => x"5997fe04",
   811 => x"a3e40880",
   812 => x"2eae387b",
   813 => x"5196e52d",
   814 => x"9ef8089e",
   815 => x"f80880ff",
   816 => x"fffff806",
   817 => x"555c7380",
   818 => x"fffffff8",
   819 => x"2e92389e",
   820 => x"f808fe05",
   821 => x"a3ec0829",
   822 => x"a3f40805",
   823 => x"5797fc04",
   824 => x"8054739e",
   825 => x"f80c02b8",
   826 => x"050d0402",
   827 => x"f4050d74",
   828 => x"70088105",
   829 => x"710c7008",
   830 => x"a3e00806",
   831 => x"5353718e",
   832 => x"38881308",
   833 => x"5196e52d",
   834 => x"9ef80888",
   835 => x"140c810b",
   836 => x"9ef80c02",
   837 => x"8c050d04",
   838 => x"02f0050d",
   839 => x"75881108",
   840 => x"fe05a3ec",
   841 => x"0829a3f4",
   842 => x"08117208",
   843 => x"a3e00806",
   844 => x"05795553",
   845 => x"54548b8c",
   846 => x"2d9ef808",
   847 => x"539ef808",
   848 => x"802e8338",
   849 => x"8153729e",
   850 => x"f80c0290",
   851 => x"050d0402",
   852 => x"ec050d77",
   853 => x"7753a3c4",
   854 => x"525397d3",
   855 => x"2d9ef808",
   856 => x"549ef808",
   857 => x"802ebf38",
   858 => x"9edc5182",
   859 => x"bb2da3c8",
   860 => x"0883ff05",
   861 => x"892a5580",
   862 => x"54737525",
   863 => x"a7387252",
   864 => x"a3c4519a",
   865 => x"982d9ef8",
   866 => x"08802e91",
   867 => x"38a3c451",
   868 => x"99eb2d84",
   869 => x"80138115",
   870 => x"55539af9",
   871 => x"049ef808",
   872 => x"549ba604",
   873 => x"8154739e",
   874 => x"f80c0294",
   875 => x"050d0400",
   876 => x"00ffffff",
   877 => x"ff00ffff",
   878 => x"ffff00ff",
   879 => x"ffffff00",
   880 => x"434d4400",
   881 => x"53504900",
   882 => x"52656164",
   883 => x"476f7420",
   884 => x"4e4f500a",
   885 => x"00000000",
   886 => x"476f7420",
   887 => x"61646472",
   888 => x"20616e64",
   889 => x"20636f75",
   890 => x"6e740a00",
   891 => x"53656e64",
   892 => x"696e6720",
   893 => x"626c6f63",
   894 => x"6b0a0000",
   895 => x"476f7420",
   896 => x"52454144",
   897 => x"43415041",
   898 => x"43495459",
   899 => x"0a000000",
   900 => x"476f7420",
   901 => x"424f4f54",
   902 => x"53545241",
   903 => x"500a0000",
   904 => x"43616e27",
   905 => x"74206f70",
   906 => x"656e2066",
   907 => x"696c650a",
   908 => x"00000000",
   909 => x"756e6b6e",
   910 => x"6f776e20",
   911 => x"636f6d6d",
   912 => x"616e640a",
   913 => x"00000000",
   914 => x"57616974",
   915 => x"696e6720",
   916 => x"666f7220",
   917 => x"6e657874",
   918 => x"20636f6d",
   919 => x"6d616e64",
   920 => x"0a000000",
   921 => x"496e6974",
   922 => x"69616c69",
   923 => x"7a696e67",
   924 => x"20534420",
   925 => x"63617264",
   926 => x"0a000000",
   927 => x"48756e74",
   928 => x"696e6720",
   929 => x"666f7220",
   930 => x"70617274",
   931 => x"6974696f",
   932 => x"6e0a0000",
   933 => x"42494f53",
   934 => x"4e455854",
   935 => x"31383600",
   936 => x"42494f53",
   937 => x"2053656e",
   938 => x"740a0000",
   939 => x"42494f53",
   940 => x"204c6f61",
   941 => x"64206661",
   942 => x"696c6564",
   943 => x"0a000000",
   944 => x"52656164",
   945 => x"696e6720",
   946 => x"4d42520a",
   947 => x"00000000",
   948 => x"52656164",
   949 => x"206f6620",
   950 => x"4d425220",
   951 => x"6661696c",
   952 => x"65640a00",
   953 => x"4d425220",
   954 => x"73756363",
   955 => x"65737366",
   956 => x"756c6c79",
   957 => x"20726561",
   958 => x"640a0000",
   959 => x"46415431",
   960 => x"36202020",
   961 => x"00000000",
   962 => x"46415433",
   963 => x"32202020",
   964 => x"00000000",
   965 => x"4e6f2070",
   966 => x"61727469",
   967 => x"74696f6e",
   968 => x"20736967",
   969 => x"6e617475",
   970 => x"72652066",
   971 => x"6f756e64",
   972 => x"0a000000",
   973 => x"52656164",
   974 => x"20626f6f",
   975 => x"74207365",
   976 => x"63746f72",
   977 => x"2066726f",
   978 => x"6d206669",
   979 => x"72737420",
   980 => x"70617274",
   981 => x"6974696f",
   982 => x"6e0a0000",
   983 => x"4f70656e",
   984 => x"65642066",
   985 => x"696c652c",
   986 => x"206c6f61",
   987 => x"64696e67",
   988 => x"2e2e2e0a",
   989 => x"002e2e0a",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba5",
     9 => x"80080b0b",
    10 => x"0ba58408",
    11 => x"0b0b0ba5",
    12 => x"88080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a5880c0b",
    16 => x"0b0ba584",
    17 => x"0c0b0b0b",
    18 => x"a5800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba2dc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a58070aa",
    57 => x"e0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8fd00402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752e80c7",
    65 => x"38875472",
    66 => x"9c2a7384",
    67 => x"2b545271",
    68 => x"802e8338",
    69 => x"81558972",
    70 => x"259938b7",
    71 => x"1252749b",
    72 => x"38ff1454",
    73 => x"738025df",
    74 => x"38800ba5",
    75 => x"800c0294",
    76 => x"050d04b0",
    77 => x"12527480",
    78 => x"2ee73871",
    79 => x"5182da2d",
    80 => x"ff145473",
    81 => x"8025c038",
    82 => x"82a904b0",
    83 => x"5182da2d",
    84 => x"800ba580",
    85 => x"0c029405",
    86 => x"0d0402f8",
    87 => x"050d7352",
    88 => x"c0087088",
    89 => x"2a708106",
    90 => x"51515170",
    91 => x"802ef138",
    92 => x"71c00c71",
    93 => x"a5800c02",
    94 => x"88050d04",
    95 => x"02f8050d",
    96 => x"7352c408",
    97 => x"70882a70",
    98 => x"81065151",
    99 => x"5170802e",
   100 => x"f13871c4",
   101 => x"0c71a580",
   102 => x"0c028805",
   103 => x"0d0402e8",
   104 => x"050d8078",
   105 => x"57557570",
   106 => x"84055708",
   107 => x"53805472",
   108 => x"982a7388",
   109 => x"2b545271",
   110 => x"802ea238",
   111 => x"c0087088",
   112 => x"2a708106",
   113 => x"51515170",
   114 => x"802ef138",
   115 => x"71c00c81",
   116 => x"15811555",
   117 => x"55837425",
   118 => x"d63871ca",
   119 => x"3874a580",
   120 => x"0c029805",
   121 => x"0d0402f4",
   122 => x"050dd452",
   123 => x"81ff720c",
   124 => x"71085381",
   125 => x"ff720c72",
   126 => x"882b83fe",
   127 => x"80067208",
   128 => x"7081ff06",
   129 => x"51525381",
   130 => x"ff720c72",
   131 => x"7107882b",
   132 => x"72087081",
   133 => x"ff065152",
   134 => x"5381ff72",
   135 => x"0c727107",
   136 => x"882b7208",
   137 => x"7081ff06",
   138 => x"7207a580",
   139 => x"0c525302",
   140 => x"8c050d04",
   141 => x"02f4050d",
   142 => x"74767181",
   143 => x"ff06d40c",
   144 => x"5353a5e4",
   145 => x"08853871",
   146 => x"892b5271",
   147 => x"982ad40c",
   148 => x"71902a70",
   149 => x"81ff06d4",
   150 => x"0c517188",
   151 => x"2a7081ff",
   152 => x"06d40c51",
   153 => x"7181ff06",
   154 => x"d40c7290",
   155 => x"2a7081ff",
   156 => x"06d40c51",
   157 => x"d4087081",
   158 => x"ff065151",
   159 => x"82b8bf52",
   160 => x"7081ff2e",
   161 => x"09810694",
   162 => x"3881ff0b",
   163 => x"d40cd408",
   164 => x"7081ff06",
   165 => x"ff145451",
   166 => x"5171e538",
   167 => x"70a5800c",
   168 => x"028c050d",
   169 => x"0402fc05",
   170 => x"0d81c751",
   171 => x"81ff0bd4",
   172 => x"0cff1151",
   173 => x"708025f4",
   174 => x"38028405",
   175 => x"0d0402f0",
   176 => x"050d85a5",
   177 => x"2d819c9f",
   178 => x"53805287",
   179 => x"fc80f751",
   180 => x"84b42da5",
   181 => x"800854a5",
   182 => x"8008812e",
   183 => x"9038ff13",
   184 => x"5372e638",
   185 => x"72a5800c",
   186 => x"0290050d",
   187 => x"0481ff0b",
   188 => x"d40c820a",
   189 => x"52849c80",
   190 => x"e95184b4",
   191 => x"2da58008",
   192 => x"802e8e38",
   193 => x"85a52dff",
   194 => x"135372ff",
   195 => x"bc3885e4",
   196 => x"0481ff0b",
   197 => x"d40c73a5",
   198 => x"800c0290",
   199 => x"050d0402",
   200 => x"f4050d81",
   201 => x"ff0bd40c",
   202 => x"a2ec5183",
   203 => x"9e2d9353",
   204 => x"805287fc",
   205 => x"80c15184",
   206 => x"b42da580",
   207 => x"08802e93",
   208 => x"3885a52d",
   209 => x"ff135372",
   210 => x"e73872a5",
   211 => x"800c028c",
   212 => x"050d0481",
   213 => x"ff0bd40c",
   214 => x"810ba580",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050d85a5",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"5184b42d",
   221 => x"a5800881",
   222 => x"2e8f3886",
   223 => x"9f2d8054",
   224 => x"73a5800c",
   225 => x"0290050d",
   226 => x"0483e62d",
   227 => x"a5800883",
   228 => x"ffff0653",
   229 => x"7283aa2e",
   230 => x"098106df",
   231 => x"3881ff0b",
   232 => x"d40cb153",
   233 => x"85be2da5",
   234 => x"80089538",
   235 => x"72822ece",
   236 => x"38ff1353",
   237 => x"72ee3872",
   238 => x"a5800c02",
   239 => x"90050d04",
   240 => x"805287fc",
   241 => x"80fa5184",
   242 => x"b42da580",
   243 => x"08de3881",
   244 => x"ff0bd40c",
   245 => x"d4085381",
   246 => x"ff0bd40c",
   247 => x"81ff0bd4",
   248 => x"0c81ff0b",
   249 => x"d40c81ff",
   250 => x"0bd40c72",
   251 => x"862a7081",
   252 => x"06a58008",
   253 => x"56515372",
   254 => x"802eff84",
   255 => x"38810ba5",
   256 => x"800c0290",
   257 => x"050d0402",
   258 => x"e8050d78",
   259 => x"5681ff0b",
   260 => x"d40cd008",
   261 => x"708f2a70",
   262 => x"81065151",
   263 => x"5372f338",
   264 => x"82810bd0",
   265 => x"0c81ff0b",
   266 => x"d40c7752",
   267 => x"87fc80d8",
   268 => x"5184b42d",
   269 => x"a5800881",
   270 => x"823881ff",
   271 => x"0bd40c81",
   272 => x"fe0bd40c",
   273 => x"80ff5575",
   274 => x"70840557",
   275 => x"0870982a",
   276 => x"d40c7090",
   277 => x"2c7081ff",
   278 => x"06d40c54",
   279 => x"70882c70",
   280 => x"81ff06d4",
   281 => x"0c547081",
   282 => x"ff06d40c",
   283 => x"54ff1555",
   284 => x"748025d3",
   285 => x"3881ff0b",
   286 => x"d40c81ff",
   287 => x"0bd40c81",
   288 => x"ff0bd40c",
   289 => x"868da054",
   290 => x"81ff0bd4",
   291 => x"0cd40881",
   292 => x"ff065574",
   293 => x"8738ff14",
   294 => x"5473ed38",
   295 => x"81ff0bd4",
   296 => x"0cd00870",
   297 => x"8f2a7081",
   298 => x"06515153",
   299 => x"72f33872",
   300 => x"d00c72a5",
   301 => x"800c0298",
   302 => x"050d04a2",
   303 => x"f051839e",
   304 => x"2d810ba5",
   305 => x"800c0298",
   306 => x"050d0402",
   307 => x"ec050d76",
   308 => x"78545480",
   309 => x"5580dbc6",
   310 => x"df5281ff",
   311 => x"0bd40cd4",
   312 => x"087081ff",
   313 => x"06515170",
   314 => x"81fe2e95",
   315 => x"38ff1252",
   316 => x"71e83881",
   317 => x"ff0bd40c",
   318 => x"74a5800c",
   319 => x"0294050d",
   320 => x"04800ba6",
   321 => x"880c8373",
   322 => x"259f3883",
   323 => x"e62da580",
   324 => x"08747084",
   325 => x"05560ca6",
   326 => x"8808a580",
   327 => x"0805a688",
   328 => x"0cfc1353",
   329 => x"728324e3",
   330 => x"38807325",
   331 => x"a03881ff",
   332 => x"0bd40cff",
   333 => x"74708105",
   334 => x"5681b72d",
   335 => x"a6880881",
   336 => x"ff05a688",
   337 => x"0cff1353",
   338 => x"728024e2",
   339 => x"38815581",
   340 => x"ff0bd40c",
   341 => x"74a5800c",
   342 => x"0294050d",
   343 => x"0402e805",
   344 => x"0d805287",
   345 => x"fc80c951",
   346 => x"84b42d92",
   347 => x"52a5f451",
   348 => x"89cb2da5",
   349 => x"f40b80f5",
   350 => x"2d81c006",
   351 => x"537280c0",
   352 => x"2e80f738",
   353 => x"a5fd0b80",
   354 => x"f52d7010",
   355 => x"8606a5fe",
   356 => x"0b80f52d",
   357 => x"70872a72",
   358 => x"07a5f90b",
   359 => x"80f52d8f",
   360 => x"06a5fa0b",
   361 => x"80f52d70",
   362 => x"8a2b9880",
   363 => x"06a5fb0b",
   364 => x"80f52d70",
   365 => x"822b7207",
   366 => x"a5fc0b80",
   367 => x"f52d7086",
   368 => x"2a720782",
   369 => x"1881782b",
   370 => x"81138173",
   371 => x"2b712951",
   372 => x"53585852",
   373 => x"52525259",
   374 => x"53545258",
   375 => x"55558480",
   376 => x"75258e38",
   377 => x"72107581",
   378 => x"2c565374",
   379 => x"848024f4",
   380 => x"3872a580",
   381 => x"0c029805",
   382 => x"0d04a5fb",
   383 => x"0b80f52d",
   384 => x"a5fc0b80",
   385 => x"f52d7190",
   386 => x"2b71882b",
   387 => x"07a5fd0b",
   388 => x"80f52d71",
   389 => x"81fffe80",
   390 => x"06077088",
   391 => x"80298880",
   392 => x"05a5800c",
   393 => x"51555755",
   394 => x"0298050d",
   395 => x"0402f405",
   396 => x"0d810ba5",
   397 => x"e40cd008",
   398 => x"708f2a70",
   399 => x"81065151",
   400 => x"5372f338",
   401 => x"72d00c85",
   402 => x"a52da380",
   403 => x"51839e2d",
   404 => x"d008708f",
   405 => x"2a708106",
   406 => x"51515372",
   407 => x"f338810b",
   408 => x"d00c8753",
   409 => x"805284d4",
   410 => x"80c05184",
   411 => x"b42da580",
   412 => x"08812e8d",
   413 => x"3872822e",
   414 => x"80c538ff",
   415 => x"135372e4",
   416 => x"3886e22d",
   417 => x"a58008a5",
   418 => x"e40ca580",
   419 => x"08802eb9",
   420 => x"3881ff0b",
   421 => x"d40c8add",
   422 => x"2da58008",
   423 => x"a5e80cd0",
   424 => x"08708f2a",
   425 => x"70810651",
   426 => x"515372f3",
   427 => x"3872d00c",
   428 => x"81ff0bd4",
   429 => x"0c810ba5",
   430 => x"800c028c",
   431 => x"050d0480",
   432 => x"0ba5800c",
   433 => x"028c050d",
   434 => x"04815287",
   435 => x"fc80d051",
   436 => x"84b42d81",
   437 => x"ff0bd40c",
   438 => x"8add2da5",
   439 => x"8008a5e8",
   440 => x"0c8d9f04",
   441 => x"02f0050d",
   442 => x"805481ff",
   443 => x"0bd40cd0",
   444 => x"08708f2a",
   445 => x"70810651",
   446 => x"515372f3",
   447 => x"3882810b",
   448 => x"d00c81ff",
   449 => x"0bd40c75",
   450 => x"5287fc80",
   451 => x"d15184b4",
   452 => x"2da58008",
   453 => x"802e8a38",
   454 => x"73a5800c",
   455 => x"0290050d",
   456 => x"04848052",
   457 => x"765189cb",
   458 => x"2da58008",
   459 => x"54d00870",
   460 => x"8f2a7081",
   461 => x"06515153",
   462 => x"72f33872",
   463 => x"d00c73a5",
   464 => x"800c0290",
   465 => x"050d0402",
   466 => x"f4050d74",
   467 => x"70882a83",
   468 => x"fe800670",
   469 => x"72982a07",
   470 => x"72882b87",
   471 => x"fc808006",
   472 => x"73982b81",
   473 => x"f00a0671",
   474 => x"730707a5",
   475 => x"800c5651",
   476 => x"5351028c",
   477 => x"050d0402",
   478 => x"f8050d02",
   479 => x"8e0580f5",
   480 => x"2d74882b",
   481 => x"077083ff",
   482 => x"ff06a580",
   483 => x"0c510288",
   484 => x"050d0402",
   485 => x"f8050d73",
   486 => x"70902b71",
   487 => x"902a07a5",
   488 => x"800c5202",
   489 => x"88050d04",
   490 => x"02f4050d",
   491 => x"a5e00853",
   492 => x"cc087082",
   493 => x"80065252",
   494 => x"70732ef4",
   495 => x"38728280",
   496 => x"32a5e00c",
   497 => x"71fdff06",
   498 => x"a5800c02",
   499 => x"8c050d04",
   500 => x"02d8050d",
   501 => x"800ba5e0",
   502 => x"0ca38451",
   503 => x"839e2d8c",
   504 => x"ad2da580",
   505 => x"088b3880",
   506 => x"0ba5800c",
   507 => x"02a8050d",
   508 => x"04a38c51",
   509 => x"839e2d97",
   510 => x"942d8fa8",
   511 => x"2da58008",
   512 => x"5aa5e008",
   513 => x"802ebc38",
   514 => x"7981822e",
   515 => x"80c53879",
   516 => x"81822482",
   517 => x"e5387984",
   518 => x"2e83c838",
   519 => x"79842485",
   520 => x"93387983",
   521 => x"2e80fb38",
   522 => x"90538052",
   523 => x"795181f7",
   524 => x"2da39451",
   525 => x"839e2d8f",
   526 => x"a82da580",
   527 => x"085aa5e0",
   528 => x"08c638a3",
   529 => x"9c51839e",
   530 => x"2d798182",
   531 => x"2e098106",
   532 => x"ffbd38a3",
   533 => x"ac51839e",
   534 => x"2da5e80b",
   535 => x"80f52da5",
   536 => x"e00807cc",
   537 => x"0c8fa82d",
   538 => x"a5e90b80",
   539 => x"f52da5e0",
   540 => x"0807cc0c",
   541 => x"8fa82da5",
   542 => x"ea0b80f5",
   543 => x"2da5e008",
   544 => x"07cc0c8f",
   545 => x"a82da5eb",
   546 => x"0b80f52d",
   547 => x"a5e00807",
   548 => x"cc0c8fa8",
   549 => x"2da58008",
   550 => x"5aa5e008",
   551 => x"feea3890",
   552 => x"c304a5e0",
   553 => x"08cc0c8f",
   554 => x"a82da580",
   555 => x"08982ba5",
   556 => x"e008cc0c",
   557 => x"588fa82d",
   558 => x"a5800890",
   559 => x"2b7807a5",
   560 => x"e008cc0c",
   561 => x"588fa82d",
   562 => x"a5800888",
   563 => x"2b7807a5",
   564 => x"e008cc0c",
   565 => x"588fa82d",
   566 => x"77a58008",
   567 => x"07a5e008",
   568 => x"cc0c588f",
   569 => x"a82da580",
   570 => x"08ff0559",
   571 => x"78ff2e80",
   572 => x"f438a6a4",
   573 => x"5779832e",
   574 => x"81bc3876",
   575 => x"52775181",
   576 => x"18588de4",
   577 => x"2d80ff56",
   578 => x"76708405",
   579 => x"58087098",
   580 => x"2aa5e008",
   581 => x"07cc0c55",
   582 => x"8fa82d74",
   583 => x"902a7081",
   584 => x"ff0670a5",
   585 => x"e00807cc",
   586 => x"0c51548f",
   587 => x"a82d7488",
   588 => x"2a7081ff",
   589 => x"0670a5e0",
   590 => x"0807cc0c",
   591 => x"51548fa8",
   592 => x"2d7481ff",
   593 => x"0670a5e0",
   594 => x"0807cc0c",
   595 => x"558fa82d",
   596 => x"ff165675",
   597 => x"8025ffb0",
   598 => x"38ff1959",
   599 => x"78ff2e09",
   600 => x"8106ff8e",
   601 => x"38a5e008",
   602 => x"cc0c8fa8",
   603 => x"2da58008",
   604 => x"5aa5e008",
   605 => x"fd923890",
   606 => x"c3047981",
   607 => x"842e80e3",
   608 => x"3881847a",
   609 => x"24fe9b38",
   610 => x"7981902e",
   611 => x"82bb3879",
   612 => x"81fe2e09",
   613 => x"8106fd90",
   614 => x"38a5e008",
   615 => x"81fe07cc",
   616 => x"0c8fa82d",
   617 => x"a5800851",
   618 => x"82da2da5",
   619 => x"e00881fe",
   620 => x"07cc0c91",
   621 => x"9204a3b4",
   622 => x"51839e2d",
   623 => x"90538052",
   624 => x"775181f7",
   625 => x"2da05182",
   626 => x"da2d7752",
   627 => x"8118aaa8",
   628 => x"5258a1a8",
   629 => x"2d7652aa",
   630 => x"a851a0ba",
   631 => x"2d80ff56",
   632 => x"928804a5",
   633 => x"e008cc0c",
   634 => x"8fa82da5",
   635 => x"8008982b",
   636 => x"a5e008cc",
   637 => x"0c588fa8",
   638 => x"2da58008",
   639 => x"902b7807",
   640 => x"a5e008cc",
   641 => x"0c588fa8",
   642 => x"2da58008",
   643 => x"882b7807",
   644 => x"a5e008cc",
   645 => x"0c588fa8",
   646 => x"2d77a580",
   647 => x"0807a5e0",
   648 => x"08cc0c58",
   649 => x"8fa82da5",
   650 => x"80085990",
   651 => x"53805277",
   652 => x"5181f72d",
   653 => x"ff195978",
   654 => x"ff2efea9",
   655 => x"38a6a40b",
   656 => x"a3b85255",
   657 => x"839e2d79",
   658 => x"842e81c8",
   659 => x"3880ff56",
   660 => x"a5e008cc",
   661 => x"0c8fa82d",
   662 => x"a5e008cc",
   663 => x"0ca58008",
   664 => x"882b548f",
   665 => x"a82da5e0",
   666 => x"08cc0c73",
   667 => x"a5800807",
   668 => x"882b548f",
   669 => x"a82da5e0",
   670 => x"08cc0c73",
   671 => x"a5800807",
   672 => x"882b548f",
   673 => x"a82d73a5",
   674 => x"80080775",
   675 => x"70840557",
   676 => x"0cff1656",
   677 => x"758025ff",
   678 => x"b738a3bc",
   679 => x"51839e2d",
   680 => x"79842e81",
   681 => x"8038a6a4",
   682 => x"52775181",
   683 => x"18588887",
   684 => x"2d94b404",
   685 => x"7981802e",
   686 => x"098106fa",
   687 => x"eb38a5e0",
   688 => x"08818007",
   689 => x"cc0c9192",
   690 => x"048056a5",
   691 => x"e008cc0c",
   692 => x"a68c1654",
   693 => x"8fa82da5",
   694 => x"80087481",
   695 => x"b72d8116",
   696 => x"568b7625",
   697 => x"e638800b",
   698 => x"a6970b81",
   699 => x"b72da68c",
   700 => x"51839e2d",
   701 => x"a68c52aa",
   702 => x"a8519dc3",
   703 => x"2da58008",
   704 => x"802eae38",
   705 => x"a5e008cc",
   706 => x"0c8fa82d",
   707 => x"a5e008cc",
   708 => x"0c92ea04",
   709 => x"77528118",
   710 => x"aaa85258",
   711 => x"a1a82d80",
   712 => x"ff5694d0",
   713 => x"04a6a452",
   714 => x"aaa851a0",
   715 => x"f12d94b4",
   716 => x"04a5e008",
   717 => x"81ff07cc",
   718 => x"0c8fa82d",
   719 => x"a5e00881",
   720 => x"ff07cc0c",
   721 => x"a3c05183",
   722 => x"9e2d90b7",
   723 => x"0402e805",
   724 => x"0d77797b",
   725 => x"58555580",
   726 => x"53727625",
   727 => x"a3387470",
   728 => x"81055680",
   729 => x"f52d7470",
   730 => x"81055680",
   731 => x"f52d5252",
   732 => x"71712e09",
   733 => x"81069338",
   734 => x"81135375",
   735 => x"7324df38",
   736 => x"800ba580",
   737 => x"0c029805",
   738 => x"0d04810b",
   739 => x"a5800c02",
   740 => x"98050d04",
   741 => x"02d8050d",
   742 => x"800baacc",
   743 => x"0ca3c851",
   744 => x"839e2da6",
   745 => x"a4528051",
   746 => x"8de42da5",
   747 => x"800854a5",
   748 => x"80089238",
   749 => x"a3d85183",
   750 => x"9e2d7356",
   751 => x"75a5800c",
   752 => x"02a8050d",
   753 => x"04a3ec51",
   754 => x"839e2d80",
   755 => x"55810ba6",
   756 => x"980c8853",
   757 => x"a48452a6",
   758 => x"da5196cd",
   759 => x"2da58008",
   760 => x"752e80fb",
   761 => x"388853a4",
   762 => x"9052a6f6",
   763 => x"5196cd2d",
   764 => x"a5800887",
   765 => x"38a58008",
   766 => x"a6980ca6",
   767 => x"9808802e",
   768 => x"818938a9",
   769 => x"ea0b80f5",
   770 => x"2da9eb0b",
   771 => x"80f52d71",
   772 => x"982b7190",
   773 => x"2b07a9ec",
   774 => x"0b80f52d",
   775 => x"70882b72",
   776 => x"07a9ed0b",
   777 => x"80f52d71",
   778 => x"07aaa20b",
   779 => x"80f52daa",
   780 => x"a30b80f5",
   781 => x"2d71882b",
   782 => x"07534055",
   783 => x"525a5657",
   784 => x"557381ab",
   785 => x"aa2ea138",
   786 => x"7382d4d5",
   787 => x"2ea338a4",
   788 => x"9c51839e",
   789 => x"2d800ba5",
   790 => x"800c02a8",
   791 => x"050d04a5",
   792 => x"8008a698",
   793 => x"0c97e504",
   794 => x"74518ec7",
   795 => x"2da58008",
   796 => x"55a6a452",
   797 => x"74518de4",
   798 => x"2da58008",
   799 => x"56a58008",
   800 => x"802efeb8",
   801 => x"38a4bc51",
   802 => x"839e2d88",
   803 => x"53a49052",
   804 => x"a6f65196",
   805 => x"cd2da580",
   806 => x"0881fa38",
   807 => x"810baacc",
   808 => x"0caaa20b",
   809 => x"80f52d54",
   810 => x"7380d52e",
   811 => x"098106ff",
   812 => x"a438aaa3",
   813 => x"0b80f52d",
   814 => x"547381aa",
   815 => x"2e098106",
   816 => x"ff933880",
   817 => x"0ba6a40b",
   818 => x"80f52d57",
   819 => x"547581e9",
   820 => x"2e833881",
   821 => x"547581eb",
   822 => x"2e8c3880",
   823 => x"5673762e",
   824 => x"098106fd",
   825 => x"d738a6af",
   826 => x"0b80f52d",
   827 => x"5675fee5",
   828 => x"38a6b00b",
   829 => x"80f52d54",
   830 => x"73822e09",
   831 => x"8106fed5",
   832 => x"38a6b10b",
   833 => x"80f52d70",
   834 => x"aad40cff",
   835 => x"05aac80c",
   836 => x"a6b20b80",
   837 => x"f52da6b3",
   838 => x"0b80f52d",
   839 => x"5b75057a",
   840 => x"82802905",
   841 => x"70aabc0c",
   842 => x"a6b40b80",
   843 => x"f52d70aa",
   844 => x"b80caacc",
   845 => x"085b5957",
   846 => x"7880f838",
   847 => x"a6b60b80",
   848 => x"f52da6b5",
   849 => x"0b80f52d",
   850 => x"71828029",
   851 => x"0570aaa4",
   852 => x"0c70a029",
   853 => x"83ff0570",
   854 => x"892a70aa",
   855 => x"d00ca6bb",
   856 => x"0b80f52d",
   857 => x"a6ba0b80",
   858 => x"f52d7182",
   859 => x"80290570",
   860 => x"a69c0c7d",
   861 => x"71291d70",
   862 => x"aac40c7f",
   863 => x"a6a00c73",
   864 => x"05aadc0c",
   865 => x"5a5a5151",
   866 => x"555a8156",
   867 => x"75a5800c",
   868 => x"02a8050d",
   869 => x"048853a4",
   870 => x"8452a6da",
   871 => x"5196cd2d",
   872 => x"8056a580",
   873 => x"08762efd",
   874 => x"f83875a5",
   875 => x"800c02a8",
   876 => x"050d0488",
   877 => x"53a49052",
   878 => x"a6f65196",
   879 => x"cd2da580",
   880 => x"08fbf938",
   881 => x"aad40870",
   882 => x"842baaa4",
   883 => x"0c70aad0",
   884 => x"0ca6c90b",
   885 => x"80f52da6",
   886 => x"c80b80f5",
   887 => x"2d718280",
   888 => x"2905a6ca",
   889 => x"0b80f52d",
   890 => x"70848080",
   891 => x"2912a6cb",
   892 => x"0b80f52d",
   893 => x"7081800a",
   894 => x"291270a6",
   895 => x"9c0caab8",
   896 => x"087129aa",
   897 => x"bc080570",
   898 => x"aadc0ca6",
   899 => x"d10b80f5",
   900 => x"2da6d00b",
   901 => x"80f52d71",
   902 => x"82802905",
   903 => x"a6d20b80",
   904 => x"f52d7084",
   905 => x"80802912",
   906 => x"a6d30b80",
   907 => x"f52d7098",
   908 => x"2b81f00a",
   909 => x"06720570",
   910 => x"a6a00cfe",
   911 => x"117e2977",
   912 => x"05aac40c",
   913 => x"52595255",
   914 => x"585e5152",
   915 => x"5f525b57",
   916 => x"55578156",
   917 => x"9b8c0402",
   918 => x"ec050d76",
   919 => x"70872c71",
   920 => x"80ff0656",
   921 => x"5653aacc",
   922 => x"088a3872",
   923 => x"882c7381",
   924 => x"ff065555",
   925 => x"a6a452aa",
   926 => x"bc081551",
   927 => x"8de42da5",
   928 => x"800853a5",
   929 => x"8008802e",
   930 => x"9c38aacc",
   931 => x"08802e9e",
   932 => x"38731010",
   933 => x"a6a40570",
   934 => x"0852538e",
   935 => x"c72da580",
   936 => x"08f00a06",
   937 => x"5372a580",
   938 => x"0c029405",
   939 => x"0d047310",
   940 => x"a6a40570",
   941 => x"80e02d52",
   942 => x"538ef72d",
   943 => x"a5800853",
   944 => x"9da50402",
   945 => x"cc050d7e",
   946 => x"605d5d80",
   947 => x"0ba6a008",
   948 => x"aac4085a",
   949 => x"5c57aacc",
   950 => x"08772e81",
   951 => x"8a38aad4",
   952 => x"08842b59",
   953 => x"80567579",
   954 => x"2780c438",
   955 => x"758f06a0",
   956 => x"18585473",
   957 => x"802e80fa",
   958 => x"38807780",
   959 => x"f52d5555",
   960 => x"73752e83",
   961 => x"38815573",
   962 => x"81e52e9a",
   963 => x"38817076",
   964 => x"06555a73",
   965 => x"802e8f38",
   966 => x"8b1780f5",
   967 => x"2d980655",
   968 => x"74802e80",
   969 => x"de388116",
   970 => x"56787626",
   971 => x"ffbe38aa",
   972 => x"cc08802e",
   973 => x"81c1387a",
   974 => x"519cd72d",
   975 => x"a58008a5",
   976 => x"800880ff",
   977 => x"fffff806",
   978 => x"555b7380",
   979 => x"fffffff8",
   980 => x"2e81a438",
   981 => x"a58008fe",
   982 => x"05aad408",
   983 => x"29aadc08",
   984 => x"05588056",
   985 => x"9de604aa",
   986 => x"d008842b",
   987 => x"5980569d",
   988 => x"e604a6a4",
   989 => x"52775181",
   990 => x"18588de4",
   991 => x"2da6a457",
   992 => x"9df9048b",
   993 => x"537b5276",
   994 => x"5196cd2d",
   995 => x"a58008ff",
   996 => x"95389c17",
   997 => x"08518ec7",
   998 => x"2da58008",
   999 => x"841e0c9a",
  1000 => x"1780e02d",
  1001 => x"518ef72d",
  1002 => x"a58008a5",
  1003 => x"80085556",
  1004 => x"aacc0897",
  1005 => x"3873881e",
  1006 => x"0c738c1e",
  1007 => x"0c747d0c",
  1008 => x"795473a5",
  1009 => x"800c02b4",
  1010 => x"050d04a5",
  1011 => x"8008881e",
  1012 => x"0c941780",
  1013 => x"e02d518e",
  1014 => x"f72da580",
  1015 => x"08902b83",
  1016 => x"fff00a06",
  1017 => x"7017707f",
  1018 => x"88050c8c",
  1019 => x"1f0c5474",
  1020 => x"7d0c7954",
  1021 => x"9fc20480",
  1022 => x"0ba5800c",
  1023 => x"02b4050d",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


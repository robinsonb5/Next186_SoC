-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba2",
     9 => x"f0080b0b",
    10 => x"0ba2f408",
    11 => x"0b0b0ba2",
    12 => x"f8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a2f80c0b",
    16 => x"0b0ba2f4",
    17 => x"0c0b0b0b",
    18 => x"a2f00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba0e4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a2f070a8",
    57 => x"d0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8efc0402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752eb538",
    65 => x"8754729c",
    66 => x"2a73842b",
    67 => x"54527180",
    68 => x"2e833881",
    69 => x"55897225",
    70 => x"8738b712",
    71 => x"5282a304",
    72 => x"b0125274",
    73 => x"802e8638",
    74 => x"715182c7",
    75 => x"2dff1454",
    76 => x"738025d2",
    77 => x"3882bd04",
    78 => x"b05182c7",
    79 => x"2d800ba2",
    80 => x"f00c0294",
    81 => x"050d0402",
    82 => x"f8050d73",
    83 => x"52c00870",
    84 => x"882a7081",
    85 => x"06515151",
    86 => x"70802ef1",
    87 => x"3871c00c",
    88 => x"71a2f00c",
    89 => x"0288050d",
    90 => x"0402f805",
    91 => x"0d7352c4",
    92 => x"0870882a",
    93 => x"70810651",
    94 => x"51517080",
    95 => x"2ef13871",
    96 => x"c40c71a2",
    97 => x"f00c0288",
    98 => x"050d0402",
    99 => x"e8050d80",
   100 => x"78575575",
   101 => x"70840557",
   102 => x"08538054",
   103 => x"72982a73",
   104 => x"882b5452",
   105 => x"71802ea2",
   106 => x"38c00870",
   107 => x"882a7081",
   108 => x"06515151",
   109 => x"70802ef1",
   110 => x"3871c00c",
   111 => x"81158115",
   112 => x"55558374",
   113 => x"25d63871",
   114 => x"ca3874a2",
   115 => x"f00c0298",
   116 => x"050d0402",
   117 => x"f4050dd4",
   118 => x"5281ff72",
   119 => x"0c710853",
   120 => x"81ff720c",
   121 => x"72882b83",
   122 => x"fe800672",
   123 => x"087081ff",
   124 => x"06515253",
   125 => x"81ff720c",
   126 => x"72710788",
   127 => x"2b720870",
   128 => x"81ff0651",
   129 => x"525381ff",
   130 => x"720c7271",
   131 => x"07882b72",
   132 => x"087081ff",
   133 => x"067207a2",
   134 => x"f00c5253",
   135 => x"028c050d",
   136 => x"0402f405",
   137 => x"0d747671",
   138 => x"81ff06d4",
   139 => x"0c5353a3",
   140 => x"d4088538",
   141 => x"71892b52",
   142 => x"71982ad4",
   143 => x"0c71902a",
   144 => x"7081ff06",
   145 => x"d40c5171",
   146 => x"882a7081",
   147 => x"ff06d40c",
   148 => x"517181ff",
   149 => x"06d40c72",
   150 => x"902a7081",
   151 => x"ff06d40c",
   152 => x"51d40870",
   153 => x"81ff0651",
   154 => x"5182b8bf",
   155 => x"527081ff",
   156 => x"2e098106",
   157 => x"943881ff",
   158 => x"0bd40cd4",
   159 => x"087081ff",
   160 => x"06ff1454",
   161 => x"515171e5",
   162 => x"3870a2f0",
   163 => x"0c028c05",
   164 => x"0d0402fc",
   165 => x"050d81c7",
   166 => x"5181ff0b",
   167 => x"d40cff11",
   168 => x"51708025",
   169 => x"f4380284",
   170 => x"050d0402",
   171 => x"f0050d85",
   172 => x"922d819c",
   173 => x"9f538052",
   174 => x"87fc80f7",
   175 => x"5184a12d",
   176 => x"a2f00854",
   177 => x"a2f00881",
   178 => x"2e098106",
   179 => x"a33881ff",
   180 => x"0bd40c82",
   181 => x"0a52849c",
   182 => x"80e95184",
   183 => x"a12da2f0",
   184 => x"088b3881",
   185 => x"ff0bd40c",
   186 => x"735385f6",
   187 => x"0485922d",
   188 => x"ff135372",
   189 => x"c13872a2",
   190 => x"f00c0290",
   191 => x"050d0402",
   192 => x"f4050d81",
   193 => x"ff0bd40c",
   194 => x"a0f45183",
   195 => x"8b2d9353",
   196 => x"805287fc",
   197 => x"80c15184",
   198 => x"a12da2f0",
   199 => x"088b3881",
   200 => x"ff0bd40c",
   201 => x"815386b2",
   202 => x"0485922d",
   203 => x"ff135372",
   204 => x"df3872a2",
   205 => x"f00c028c",
   206 => x"050d0402",
   207 => x"f0050d85",
   208 => x"922d83aa",
   209 => x"52849c80",
   210 => x"c85184a1",
   211 => x"2da2f008",
   212 => x"812e0981",
   213 => x"06923883",
   214 => x"d32da2f0",
   215 => x"0883ffff",
   216 => x"06537283",
   217 => x"aa2e9138",
   218 => x"85ff2d86",
   219 => x"f3048154",
   220 => x"87d80480",
   221 => x"5487d804",
   222 => x"81ff0bd4",
   223 => x"0cb15385",
   224 => x"ab2da2f0",
   225 => x"08802e80",
   226 => x"c0388052",
   227 => x"87fc80fa",
   228 => x"5184a12d",
   229 => x"a2f008b1",
   230 => x"3881ff0b",
   231 => x"d40cd408",
   232 => x"5381ff0b",
   233 => x"d40c81ff",
   234 => x"0bd40c81",
   235 => x"ff0bd40c",
   236 => x"81ff0bd4",
   237 => x"0c72862a",
   238 => x"708106a2",
   239 => x"f0085651",
   240 => x"5372802e",
   241 => x"933886ee",
   242 => x"0472822e",
   243 => x"ffa538ff",
   244 => x"135372ff",
   245 => x"aa387254",
   246 => x"73a2f00c",
   247 => x"0290050d",
   248 => x"0402e805",
   249 => x"0d785681",
   250 => x"ff0bd40c",
   251 => x"d008708f",
   252 => x"2a708106",
   253 => x"51515372",
   254 => x"f3388281",
   255 => x"0bd00c81",
   256 => x"ff0bd40c",
   257 => x"775287fc",
   258 => x"80d85184",
   259 => x"a12da2f0",
   260 => x"08802e8c",
   261 => x"38a0f851",
   262 => x"838b2d81",
   263 => x"53899804",
   264 => x"81ff0bd4",
   265 => x"0c81fe0b",
   266 => x"d40c80ff",
   267 => x"55757084",
   268 => x"05570870",
   269 => x"982ad40c",
   270 => x"70902c70",
   271 => x"81ff06d4",
   272 => x"0c547088",
   273 => x"2c7081ff",
   274 => x"06d40c54",
   275 => x"7081ff06",
   276 => x"d40c54ff",
   277 => x"15557480",
   278 => x"25d33881",
   279 => x"ff0bd40c",
   280 => x"81ff0bd4",
   281 => x"0c81ff0b",
   282 => x"d40c868d",
   283 => x"a05481ff",
   284 => x"0bd40cd4",
   285 => x"0881ff06",
   286 => x"55748738",
   287 => x"ff145473",
   288 => x"ed3881ff",
   289 => x"0bd40cd0",
   290 => x"08708f2a",
   291 => x"70810651",
   292 => x"515372f3",
   293 => x"3872d00c",
   294 => x"72a2f00c",
   295 => x"0298050d",
   296 => x"0402ec05",
   297 => x"0d767853",
   298 => x"54805580",
   299 => x"dbc6df53",
   300 => x"81ff0bd4",
   301 => x"0cd40870",
   302 => x"81ff0651",
   303 => x"517081fe",
   304 => x"2e098106",
   305 => x"80ce3880",
   306 => x"0ba3f80c",
   307 => x"8372259d",
   308 => x"3883d32d",
   309 => x"a2f00874",
   310 => x"70840556",
   311 => x"0ca3f808",
   312 => x"a2f00805",
   313 => x"a3f80cfc",
   314 => x"125289cc",
   315 => x"04807225",
   316 => x"9e3881ff",
   317 => x"0bd40cff",
   318 => x"74708105",
   319 => x"5681b72d",
   320 => x"a3f80881",
   321 => x"ff05a3f8",
   322 => x"0cff1252",
   323 => x"89ed0481",
   324 => x"558a9b04",
   325 => x"ff135372",
   326 => x"ff963881",
   327 => x"ff0bd40c",
   328 => x"74a2f00c",
   329 => x"0294050d",
   330 => x"0402e805",
   331 => x"0d805287",
   332 => x"fc80c951",
   333 => x"84a12d92",
   334 => x"52a3e451",
   335 => x"89a12da3",
   336 => x"e40b80f5",
   337 => x"2d81c006",
   338 => x"537280c0",
   339 => x"2e098106",
   340 => x"b038a3eb",
   341 => x"0b80f52d",
   342 => x"a3ec0b80",
   343 => x"f52d7190",
   344 => x"2b71882b",
   345 => x"07a3ed0b",
   346 => x"80f52d71",
   347 => x"81fffe80",
   348 => x"06077088",
   349 => x"80298880",
   350 => x"05515155",
   351 => x"57558beb",
   352 => x"04a3ed0b",
   353 => x"80f52d70",
   354 => x"108606a3",
   355 => x"ee0b80f5",
   356 => x"2d70872a",
   357 => x"7207a3e9",
   358 => x"0b80f52d",
   359 => x"8f06a3ea",
   360 => x"0b80f52d",
   361 => x"708a2b98",
   362 => x"8006a3eb",
   363 => x"0b80f52d",
   364 => x"70822b72",
   365 => x"07a3ec0b",
   366 => x"80f52d70",
   367 => x"862a7207",
   368 => x"82188178",
   369 => x"2b811381",
   370 => x"732b7129",
   371 => x"51535858",
   372 => x"52525252",
   373 => x"59535452",
   374 => x"58555584",
   375 => x"8075258b",
   376 => x"38721075",
   377 => x"812c5653",
   378 => x"8bdb0472",
   379 => x"a2f00c02",
   380 => x"98050d04",
   381 => x"02f0050d",
   382 => x"810ba3d4",
   383 => x"0ca18851",
   384 => x"838b2d87",
   385 => x"54d00870",
   386 => x"8f2a7081",
   387 => x"06515153",
   388 => x"72f33872",
   389 => x"d00c8592",
   390 => x"2dd00870",
   391 => x"8f2a7081",
   392 => x"06515153",
   393 => x"72f33881",
   394 => x"0bd00c72",
   395 => x"5284d480",
   396 => x"c05184a1",
   397 => x"2da2f008",
   398 => x"812e9938",
   399 => x"73822e09",
   400 => x"81068a38",
   401 => x"a18c5183",
   402 => x"8b2d8d92",
   403 => x"04ff1454",
   404 => x"73ffb238",
   405 => x"86bb2da2",
   406 => x"f008a3d4",
   407 => x"0ca2f008",
   408 => x"8b388152",
   409 => x"87fc80d0",
   410 => x"5184a12d",
   411 => x"81ff0bd4",
   412 => x"0c8aa92d",
   413 => x"a2f008a3",
   414 => x"d80cd008",
   415 => x"708f2a70",
   416 => x"81065151",
   417 => x"5372f338",
   418 => x"72d00c81",
   419 => x"ff0bd40c",
   420 => x"815372a2",
   421 => x"f00c0290",
   422 => x"050d0402",
   423 => x"f0050d80",
   424 => x"5481ff0b",
   425 => x"d40cd008",
   426 => x"708f2a70",
   427 => x"81065151",
   428 => x"5372f338",
   429 => x"82810bd0",
   430 => x"0c81ff0b",
   431 => x"d40c7552",
   432 => x"87fc80d1",
   433 => x"5184a12d",
   434 => x"a2f0089e",
   435 => x"38848052",
   436 => x"765189a1",
   437 => x"2da2f008",
   438 => x"54d00870",
   439 => x"8f2a7081",
   440 => x"06515153",
   441 => x"72f33872",
   442 => x"d00c73a2",
   443 => x"f00c0290",
   444 => x"050d0402",
   445 => x"f4050d74",
   446 => x"70882a83",
   447 => x"fe800670",
   448 => x"72982a07",
   449 => x"72882b87",
   450 => x"fc808006",
   451 => x"73982b81",
   452 => x"f00a0671",
   453 => x"730707a2",
   454 => x"f00c5651",
   455 => x"5351028c",
   456 => x"050d0402",
   457 => x"f8050d02",
   458 => x"8e0580f5",
   459 => x"2d74882b",
   460 => x"077083ff",
   461 => x"ff06a2f0",
   462 => x"0c510288",
   463 => x"050d0402",
   464 => x"f8050d73",
   465 => x"70902b71",
   466 => x"902a07a2",
   467 => x"f00c5202",
   468 => x"88050d04",
   469 => x"02f4050d",
   470 => x"a3d00853",
   471 => x"cc087082",
   472 => x"80065252",
   473 => x"70732ef4",
   474 => x"38728280",
   475 => x"32a3d00c",
   476 => x"71fdff06",
   477 => x"a2f00c02",
   478 => x"8c050d04",
   479 => x"02d8050d",
   480 => x"800ba3d0",
   481 => x"0ca19451",
   482 => x"838b2d8b",
   483 => x"f42da2f0",
   484 => x"08802e86",
   485 => x"8f38a19c",
   486 => x"51838b2d",
   487 => x"95ec2d8e",
   488 => x"d42da2f0",
   489 => x"085aa2f0",
   490 => x"0881822e",
   491 => x"85a038a2",
   492 => x"f0088182",
   493 => x"24a638a2",
   494 => x"f008842e",
   495 => x"81ca38a2",
   496 => x"f0088424",
   497 => x"8c38a2f0",
   498 => x"08832e83",
   499 => x"97389592",
   500 => x"04a2f008",
   501 => x"81802eab",
   502 => x"38959204",
   503 => x"a2f00881",
   504 => x"842e81a4",
   505 => x"3881840b",
   506 => x"a2f00824",
   507 => x"82f638a2",
   508 => x"f0088190",
   509 => x"2e9738a2",
   510 => x"f00881fe",
   511 => x"2e80ed38",
   512 => x"959204a3",
   513 => x"d0088180",
   514 => x"0754958c",
   515 => x"048058a3",
   516 => x"d008cc0c",
   517 => x"a3fc1854",
   518 => x"8ed42da2",
   519 => x"f0087481",
   520 => x"b72d8118",
   521 => x"588b7825",
   522 => x"e638800b",
   523 => x"a4870b81",
   524 => x"b72da3fc",
   525 => x"51838b2d",
   526 => x"a3fc52a8",
   527 => x"98519c90",
   528 => x"2da2f008",
   529 => x"802e8c38",
   530 => x"a3d008cc",
   531 => x"0c8ed42d",
   532 => x"94c604a3",
   533 => x"d00881ff",
   534 => x"07cc0c8e",
   535 => x"d42da3d0",
   536 => x"0881ff07",
   537 => x"cc0ca1a4",
   538 => x"51959e04",
   539 => x"a3d00881",
   540 => x"fe07cc0c",
   541 => x"8ed42da2",
   542 => x"f0085182",
   543 => x"c72da3d0",
   544 => x"0881fe07",
   545 => x"54958c04",
   546 => x"a3d008cc",
   547 => x"0c8ed42d",
   548 => x"a2f00898",
   549 => x"2ba3d008",
   550 => x"cc0c568e",
   551 => x"d42da2f0",
   552 => x"08902b76",
   553 => x"07a3d008",
   554 => x"cc0c568e",
   555 => x"d42da2f0",
   556 => x"08882b76",
   557 => x"07a3d008",
   558 => x"cc0c568e",
   559 => x"d42d75a2",
   560 => x"f00807a3",
   561 => x"d008cc0c",
   562 => x"568ed42d",
   563 => x"a2f00857",
   564 => x"80f75182",
   565 => x"c72dff17",
   566 => x"5776ff2e",
   567 => x"82e838a4",
   568 => x"94557984",
   569 => x"2e098106",
   570 => x"8c387552",
   571 => x"8116a898",
   572 => x"52569fc7",
   573 => x"2d80ff58",
   574 => x"a3d008cc",
   575 => x"0c8ed42d",
   576 => x"a3d008cc",
   577 => x"0ca2f008",
   578 => x"882b548e",
   579 => x"d42da3d0",
   580 => x"08cc0c73",
   581 => x"a2f00807",
   582 => x"882b548e",
   583 => x"d42da3d0",
   584 => x"08cc0c73",
   585 => x"a2f00807",
   586 => x"882b548e",
   587 => x"d42d73a2",
   588 => x"f0080775",
   589 => x"70840557",
   590 => x"0cff1858",
   591 => x"778025ff",
   592 => x"b7387984",
   593 => x"2e098106",
   594 => x"8d38a494",
   595 => x"52a89851",
   596 => x"9f902d91",
   597 => x"d604a494",
   598 => x"52755181",
   599 => x"165687e1",
   600 => x"2d91d604",
   601 => x"80f25182",
   602 => x"c72da3d0",
   603 => x"08cc0c8e",
   604 => x"d42da2f0",
   605 => x"08982ba3",
   606 => x"d008cc0c",
   607 => x"568ed42d",
   608 => x"a2f00890",
   609 => x"2b7607a3",
   610 => x"d008cc0c",
   611 => x"568ed42d",
   612 => x"a2f00888",
   613 => x"2b7607a3",
   614 => x"d008cc0c",
   615 => x"568ed42d",
   616 => x"75a2f008",
   617 => x"07a3d008",
   618 => x"cc0c568e",
   619 => x"d42da2f0",
   620 => x"08ff0557",
   621 => x"76ff2e81",
   622 => x"8d38a494",
   623 => x"0b811755",
   624 => x"5979832e",
   625 => x"0981069b",
   626 => x"38a05182",
   627 => x"c72d7552",
   628 => x"73a89852",
   629 => x"569fc72d",
   630 => x"7852a898",
   631 => x"519ed92d",
   632 => x"93ec0478",
   633 => x"52755173",
   634 => x"568d9b2d",
   635 => x"80ff5878",
   636 => x"7084055a",
   637 => x"0870982a",
   638 => x"a3d00807",
   639 => x"cc0c558e",
   640 => x"d42d7490",
   641 => x"2a7081ff",
   642 => x"0670a3d0",
   643 => x"0807cc0c",
   644 => x"51548ed4",
   645 => x"2d74882a",
   646 => x"7081ff06",
   647 => x"70a3d008",
   648 => x"07cc0c51",
   649 => x"548ed42d",
   650 => x"7481ff06",
   651 => x"70a3d008",
   652 => x"07cc0c55",
   653 => x"8ed42dff",
   654 => x"18587780",
   655 => x"25ffb038",
   656 => x"ff175793",
   657 => x"b404a3d0",
   658 => x"08cc0c8f",
   659 => x"9f04a1ac",
   660 => x"51838b2d",
   661 => x"a3d80b80",
   662 => x"f52da3d0",
   663 => x"0807cc0c",
   664 => x"8ed42da3",
   665 => x"d90b80f5",
   666 => x"2da3d008",
   667 => x"07cc0c8e",
   668 => x"d42da3da",
   669 => x"0b80f52d",
   670 => x"a3d00807",
   671 => x"cc0c8ed4",
   672 => x"2da3db0b",
   673 => x"80f52da3",
   674 => x"d0080754",
   675 => x"73cc0c8f",
   676 => x"9f049053",
   677 => x"80527951",
   678 => x"81f72da1",
   679 => x"b451838b",
   680 => x"2d8f9f04",
   681 => x"800ba2f0",
   682 => x"0c02a805",
   683 => x"0d0402e8",
   684 => x"050d7779",
   685 => x"7b585555",
   686 => x"80537276",
   687 => x"25a33874",
   688 => x"70810556",
   689 => x"80f52d74",
   690 => x"70810556",
   691 => x"80f52d52",
   692 => x"5271712e",
   693 => x"86388151",
   694 => x"95e30481",
   695 => x"135395ba",
   696 => x"04805170",
   697 => x"a2f00c02",
   698 => x"98050d04",
   699 => x"02d8050d",
   700 => x"800ba8bc",
   701 => x"0ca1b851",
   702 => x"838b2da4",
   703 => x"94528051",
   704 => x"8d9b2da2",
   705 => x"f00854a2",
   706 => x"f0088c38",
   707 => x"a1c85183",
   708 => x"8b2d7355",
   709 => x"9b9904a1",
   710 => x"dc51838b",
   711 => x"2d805681",
   712 => x"0ba4880c",
   713 => x"8853a1f4",
   714 => x"52a4ca51",
   715 => x"95ae2da2",
   716 => x"f008762e",
   717 => x"09810687",
   718 => x"38a2f008",
   719 => x"a4880c88",
   720 => x"53a28052",
   721 => x"a4e65195",
   722 => x"ae2da2f0",
   723 => x"088738a2",
   724 => x"f008a488",
   725 => x"0ca48808",
   726 => x"802e80ff",
   727 => x"38a7da0b",
   728 => x"80f52da7",
   729 => x"db0b80f5",
   730 => x"2d71982b",
   731 => x"71902b07",
   732 => x"a7dc0b80",
   733 => x"f52d7088",
   734 => x"2b7207a7",
   735 => x"dd0b80f5",
   736 => x"2d7107a8",
   737 => x"920b80f5",
   738 => x"2da8930b",
   739 => x"80f52d71",
   740 => x"882b0753",
   741 => x"5f54525a",
   742 => x"56575573",
   743 => x"81abaa2e",
   744 => x"0981068d",
   745 => x"3875518d",
   746 => x"f32da2f0",
   747 => x"085697c1",
   748 => x"047382d4",
   749 => x"d52e8a38",
   750 => x"a28c5183",
   751 => x"8b2d98e5",
   752 => x"04a49452",
   753 => x"75518d9b",
   754 => x"2da2f008",
   755 => x"55a2f008",
   756 => x"802e83c5",
   757 => x"38a2ac51",
   758 => x"838b2d88",
   759 => x"53a28052",
   760 => x"a4e65195",
   761 => x"ae2da2f0",
   762 => x"08893881",
   763 => x"0ba8bc0c",
   764 => x"988b0488",
   765 => x"53a1f452",
   766 => x"a4ca5195",
   767 => x"ae2d8055",
   768 => x"a2f00875",
   769 => x"2e098106",
   770 => x"838f38a8",
   771 => x"920b80f5",
   772 => x"2d547380",
   773 => x"d52e0981",
   774 => x"0680ca38",
   775 => x"a8930b80",
   776 => x"f52d5473",
   777 => x"81aa2e09",
   778 => x"8106ba38",
   779 => x"800ba494",
   780 => x"0b80f52d",
   781 => x"56547481",
   782 => x"e92e8338",
   783 => x"81547481",
   784 => x"eb2e8c38",
   785 => x"80557375",
   786 => x"2e098106",
   787 => x"82cb38a4",
   788 => x"9f0b80f5",
   789 => x"2d55748d",
   790 => x"38a4a00b",
   791 => x"80f52d54",
   792 => x"73822e86",
   793 => x"3880559b",
   794 => x"9904a4a1",
   795 => x"0b80f52d",
   796 => x"70a8c40c",
   797 => x"ff05a8b8",
   798 => x"0ca4a20b",
   799 => x"80f52da4",
   800 => x"a30b80f5",
   801 => x"2d587605",
   802 => x"77828029",
   803 => x"0570a8ac",
   804 => x"0ca4a40b",
   805 => x"80f52d70",
   806 => x"a8a80ca8",
   807 => x"bc085957",
   808 => x"5876802e",
   809 => x"81a33888",
   810 => x"53a28052",
   811 => x"a4e65195",
   812 => x"ae2da2f0",
   813 => x"0881e238",
   814 => x"a8c40870",
   815 => x"842ba894",
   816 => x"0c70a8c0",
   817 => x"0ca4b90b",
   818 => x"80f52da4",
   819 => x"b80b80f5",
   820 => x"2d718280",
   821 => x"2905a4ba",
   822 => x"0b80f52d",
   823 => x"70848080",
   824 => x"2912a4bb",
   825 => x"0b80f52d",
   826 => x"7081800a",
   827 => x"291270a4",
   828 => x"8c0ca8a8",
   829 => x"087129a8",
   830 => x"ac080570",
   831 => x"a8cc0ca4",
   832 => x"c10b80f5",
   833 => x"2da4c00b",
   834 => x"80f52d71",
   835 => x"82802905",
   836 => x"a4c20b80",
   837 => x"f52d7084",
   838 => x"80802912",
   839 => x"a4c30b80",
   840 => x"f52d7098",
   841 => x"2b81f00a",
   842 => x"06720570",
   843 => x"a4900cfe",
   844 => x"117e2977",
   845 => x"05a8b40c",
   846 => x"52595243",
   847 => x"545e5152",
   848 => x"59525d57",
   849 => x"59579b97",
   850 => x"04a4a60b",
   851 => x"80f52da4",
   852 => x"a50b80f5",
   853 => x"2d718280",
   854 => x"290570a8",
   855 => x"940c70a0",
   856 => x"2983ff05",
   857 => x"70892a70",
   858 => x"a8c00ca4",
   859 => x"ab0b80f5",
   860 => x"2da4aa0b",
   861 => x"80f52d71",
   862 => x"82802905",
   863 => x"70a48c0c",
   864 => x"7b71291e",
   865 => x"70a8b40c",
   866 => x"7da4900c",
   867 => x"7305a8cc",
   868 => x"0c555e51",
   869 => x"51555581",
   870 => x"5574a2f0",
   871 => x"0c02a805",
   872 => x"0d0402ec",
   873 => x"050d7670",
   874 => x"872c7180",
   875 => x"ff065556",
   876 => x"54a8bc08",
   877 => x"8a387388",
   878 => x"2c7481ff",
   879 => x"065455a4",
   880 => x"9452a8ac",
   881 => x"0815518d",
   882 => x"9b2da2f0",
   883 => x"0854a2f0",
   884 => x"08802eb3",
   885 => x"38a8bc08",
   886 => x"802e9838",
   887 => x"728429a4",
   888 => x"94057008",
   889 => x"52538df3",
   890 => x"2da2f008",
   891 => x"f00a0653",
   892 => x"9c850472",
   893 => x"10a49405",
   894 => x"7080e02d",
   895 => x"52538ea3",
   896 => x"2da2f008",
   897 => x"53725473",
   898 => x"a2f00c02",
   899 => x"94050d04",
   900 => x"02c8050d",
   901 => x"7f615f5b",
   902 => x"800ba490",
   903 => x"08a8b408",
   904 => x"595d56a8",
   905 => x"bc08762e",
   906 => x"8a38a8c4",
   907 => x"08842b58",
   908 => x"9cb904a8",
   909 => x"c008842b",
   910 => x"58805978",
   911 => x"782781ad",
   912 => x"38788f06",
   913 => x"a0175754",
   914 => x"738f38a4",
   915 => x"94527651",
   916 => x"8117578d",
   917 => x"9b2da494",
   918 => x"56807680",
   919 => x"f52d5654",
   920 => x"74742e83",
   921 => x"38815474",
   922 => x"81e52e80",
   923 => x"fa388170",
   924 => x"7506555d",
   925 => x"73802e80",
   926 => x"ee388b16",
   927 => x"80f52d98",
   928 => x"065a7980",
   929 => x"e2388b53",
   930 => x"7d527551",
   931 => x"95ae2da2",
   932 => x"f00880d3",
   933 => x"389c1608",
   934 => x"518df32d",
   935 => x"a2f00884",
   936 => x"1c0c9a16",
   937 => x"80e02d51",
   938 => x"8ea32da2",
   939 => x"f008a2f0",
   940 => x"08881d0c",
   941 => x"a2f00855",
   942 => x"55a8bc08",
   943 => x"802e9838",
   944 => x"941680e0",
   945 => x"2d518ea3",
   946 => x"2da2f008",
   947 => x"902b83ff",
   948 => x"f00a0670",
   949 => x"16515473",
   950 => x"881c0c73",
   951 => x"8c1c0c79",
   952 => x"7b0c7c54",
   953 => x"9ea30481",
   954 => x"19599cbb",
   955 => x"04a8bc08",
   956 => x"802eae38",
   957 => x"7b519ba2",
   958 => x"2da2f008",
   959 => x"a2f00880",
   960 => x"fffffff8",
   961 => x"06555c73",
   962 => x"80ffffff",
   963 => x"f82e9238",
   964 => x"a2f008fe",
   965 => x"05a8c408",
   966 => x"29a8cc08",
   967 => x"05579cb9",
   968 => x"04805473",
   969 => x"a2f00c02",
   970 => x"b8050d04",
   971 => x"02f4050d",
   972 => x"74700881",
   973 => x"05710c70",
   974 => x"08a8b808",
   975 => x"06535371",
   976 => x"8e388813",
   977 => x"08519ba2",
   978 => x"2da2f008",
   979 => x"88140c81",
   980 => x"0ba2f00c",
   981 => x"028c050d",
   982 => x"0402f005",
   983 => x"0d758811",
   984 => x"08fe05a8",
   985 => x"c40829a8",
   986 => x"cc081172",
   987 => x"08a8b808",
   988 => x"06057955",
   989 => x"5354548d",
   990 => x"9b2da2f0",
   991 => x"0853a2f0",
   992 => x"08802e83",
   993 => x"38815372",
   994 => x"a2f00c02",
   995 => x"90050d04",
   996 => x"02f0050d",
   997 => x"75881108",
   998 => x"fe05a8c4",
   999 => x"0829a8cc",
  1000 => x"08117208",
  1001 => x"a8b80806",
  1002 => x"05795553",
  1003 => x"545487e1",
  1004 => x"2da2f008",
  1005 => x"53a2f008",
  1006 => x"802e8338",
  1007 => x"815372a2",
  1008 => x"f00c0290",
  1009 => x"050d0402",
  1010 => x"ec050d76",
  1011 => x"78841208",
  1012 => x"892a5455",
  1013 => x"53805573",
  1014 => x"7227a038",
  1015 => x"73730827",
  1016 => x"8a387473",
  1017 => x"0c8c1308",
  1018 => x"88140c72",
  1019 => x"08742e89",
  1020 => x"3872519e",
  1021 => x"ac2d9feb",
  1022 => x"04815574",
  1023 => x"a2f00c02",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


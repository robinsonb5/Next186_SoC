-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0b9c",
     9 => x"e4080b0b",
    10 => x"0b9ce808",
    11 => x"0b0b0b9c",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"9cec0c0b",
    16 => x"0b0b9ce8",
    17 => x"0c0b0b0b",
    18 => x"9ce40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b99d8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"9ce470a1",
    57 => x"e4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8ed80402",
    62 => x"f8050d73",
    63 => x"52c00870",
    64 => x"882a7081",
    65 => x"06515151",
    66 => x"70802ef1",
    67 => x"3871c00c",
    68 => x"719ce40c",
    69 => x"0288050d",
    70 => x"0402f805",
    71 => x"0d7352c4",
    72 => x"0870882a",
    73 => x"70810651",
    74 => x"51517080",
    75 => x"2ef13871",
    76 => x"c40c719c",
    77 => x"e40c0288",
    78 => x"050d0402",
    79 => x"e8050d80",
    80 => x"78575575",
    81 => x"70840557",
    82 => x"08538054",
    83 => x"72982a73",
    84 => x"882b5452",
    85 => x"71802ea2",
    86 => x"38c00870",
    87 => x"882a7081",
    88 => x"06515151",
    89 => x"70802ef1",
    90 => x"3871c00c",
    91 => x"81158115",
    92 => x"55558374",
    93 => x"25d63871",
    94 => x"ca38749c",
    95 => x"e40c0298",
    96 => x"050d0402",
    97 => x"f8050dc0",
    98 => x"0870892a",
    99 => x"70810651",
   100 => x"52527080",
   101 => x"2ef13871",
   102 => x"81ff069c",
   103 => x"e40c0288",
   104 => x"050d0402",
   105 => x"f4050dd4",
   106 => x"5281ff72",
   107 => x"0c710853",
   108 => x"81ff720c",
   109 => x"72882b83",
   110 => x"fe800672",
   111 => x"087081ff",
   112 => x"06515253",
   113 => x"81ff720c",
   114 => x"72710788",
   115 => x"2b720870",
   116 => x"81ff0651",
   117 => x"525381ff",
   118 => x"720c7271",
   119 => x"07882b72",
   120 => x"087081ff",
   121 => x"0672079c",
   122 => x"e40c5253",
   123 => x"028c050d",
   124 => x"0402f405",
   125 => x"0d747671",
   126 => x"81ff06d4",
   127 => x"0c53539c",
   128 => x"f8088538",
   129 => x"71892b52",
   130 => x"71982ad4",
   131 => x"0c71902a",
   132 => x"7081ff06",
   133 => x"d40c5171",
   134 => x"882a7081",
   135 => x"ff06d40c",
   136 => x"517181ff",
   137 => x"06d40c72",
   138 => x"902a7081",
   139 => x"ff06d40c",
   140 => x"51d40870",
   141 => x"81ff0651",
   142 => x"5182b8bf",
   143 => x"527081ff",
   144 => x"2e098106",
   145 => x"943881ff",
   146 => x"0bd40cd4",
   147 => x"087081ff",
   148 => x"06ff1454",
   149 => x"515171e5",
   150 => x"38709ce4",
   151 => x"0c028c05",
   152 => x"0d0402fc",
   153 => x"050d81c7",
   154 => x"5181ff0b",
   155 => x"d40cff11",
   156 => x"51708025",
   157 => x"f4380284",
   158 => x"050d0402",
   159 => x"f0050d84",
   160 => x"e22d819c",
   161 => x"9f538052",
   162 => x"87fc80f7",
   163 => x"5183f12d",
   164 => x"9ce40854",
   165 => x"9ce40881",
   166 => x"2e098106",
   167 => x"a33881ff",
   168 => x"0bd40c82",
   169 => x"0a52849c",
   170 => x"80e95183",
   171 => x"f12d9ce4",
   172 => x"088b3881",
   173 => x"ff0bd40c",
   174 => x"735385c6",
   175 => x"0484e22d",
   176 => x"ff135372",
   177 => x"c138729c",
   178 => x"e40c0290",
   179 => x"050d0402",
   180 => x"f4050d81",
   181 => x"ff0bd40c",
   182 => x"99e85182",
   183 => x"bb2d9353",
   184 => x"805287fc",
   185 => x"80c15183",
   186 => x"f12d9ce4",
   187 => x"088b3881",
   188 => x"ff0bd40c",
   189 => x"81538682",
   190 => x"0484e22d",
   191 => x"ff135372",
   192 => x"df38729c",
   193 => x"e40c028c",
   194 => x"050d0402",
   195 => x"f0050d84",
   196 => x"e22d83aa",
   197 => x"52849c80",
   198 => x"c85183f1",
   199 => x"2d9ce408",
   200 => x"812e0981",
   201 => x"06923883",
   202 => x"a32d9ce4",
   203 => x"0883ffff",
   204 => x"06537283",
   205 => x"aa2e9138",
   206 => x"85cf2d86",
   207 => x"c3048154",
   208 => x"87a80480",
   209 => x"5487a804",
   210 => x"81ff0bd4",
   211 => x"0cb15384",
   212 => x"fb2d9ce4",
   213 => x"08802e80",
   214 => x"c0388052",
   215 => x"87fc80fa",
   216 => x"5183f12d",
   217 => x"9ce408b1",
   218 => x"3881ff0b",
   219 => x"d40cd408",
   220 => x"5381ff0b",
   221 => x"d40c81ff",
   222 => x"0bd40c81",
   223 => x"ff0bd40c",
   224 => x"81ff0bd4",
   225 => x"0c72862a",
   226 => x"7081069c",
   227 => x"e4085651",
   228 => x"5372802e",
   229 => x"933886be",
   230 => x"0472822e",
   231 => x"ffa538ff",
   232 => x"135372ff",
   233 => x"aa387254",
   234 => x"739ce40c",
   235 => x"0290050d",
   236 => x"04800b9c",
   237 => x"e40c0402",
   238 => x"ec050d76",
   239 => x"78535480",
   240 => x"5580dbc6",
   241 => x"df5381ff",
   242 => x"0bd40cd4",
   243 => x"087081ff",
   244 => x"06515170",
   245 => x"81fe2e09",
   246 => x"810680ce",
   247 => x"38800b9d",
   248 => x"9c0c8372",
   249 => x"259d3883",
   250 => x"a32d9ce4",
   251 => x"08747084",
   252 => x"05560c9d",
   253 => x"9c089ce4",
   254 => x"08059d9c",
   255 => x"0cfc1252",
   256 => x"87e20480",
   257 => x"72259e38",
   258 => x"81ff0bd4",
   259 => x"0cff7470",
   260 => x"81055681",
   261 => x"b72d9d9c",
   262 => x"0881ff05",
   263 => x"9d9c0cff",
   264 => x"12528883",
   265 => x"04815588",
   266 => x"b104ff13",
   267 => x"5372ff96",
   268 => x"3881ff0b",
   269 => x"d40c749c",
   270 => x"e40c0294",
   271 => x"050d0402",
   272 => x"e8050d80",
   273 => x"5287fc80",
   274 => x"c95183f1",
   275 => x"2d92529d",
   276 => x"885187b7",
   277 => x"2d9d880b",
   278 => x"80f52d81",
   279 => x"c0065372",
   280 => x"80c02e09",
   281 => x"8106b038",
   282 => x"9d8f0b80",
   283 => x"f52d9d90",
   284 => x"0b80f52d",
   285 => x"71902b71",
   286 => x"882b079d",
   287 => x"910b80f5",
   288 => x"2d7181ff",
   289 => x"fe800607",
   290 => x"70888029",
   291 => x"88800551",
   292 => x"51555755",
   293 => x"8a81049d",
   294 => x"910b80f5",
   295 => x"2d701086",
   296 => x"069d920b",
   297 => x"80f52d70",
   298 => x"872a7207",
   299 => x"9d8d0b80",
   300 => x"f52d8f06",
   301 => x"9d8e0b80",
   302 => x"f52d708a",
   303 => x"2b988006",
   304 => x"9d8f0b80",
   305 => x"f52d7082",
   306 => x"2b72079d",
   307 => x"900b80f5",
   308 => x"2d70862a",
   309 => x"72078218",
   310 => x"81782b81",
   311 => x"1381732b",
   312 => x"71295153",
   313 => x"58585252",
   314 => x"52525953",
   315 => x"54525855",
   316 => x"55848075",
   317 => x"258b3872",
   318 => x"1075812c",
   319 => x"565389f1",
   320 => x"04729ce4",
   321 => x"0c029805",
   322 => x"0d0402f4",
   323 => x"050d810b",
   324 => x"9cf80cd0",
   325 => x"08708f2a",
   326 => x"70810651",
   327 => x"515372f3",
   328 => x"3872d00c",
   329 => x"84e22d99",
   330 => x"ec5182bb",
   331 => x"2dd00870",
   332 => x"8f2a7081",
   333 => x"06515153",
   334 => x"72f33881",
   335 => x"0bd00c87",
   336 => x"53805284",
   337 => x"d480c051",
   338 => x"83f12d9c",
   339 => x"e408812e",
   340 => x"94387282",
   341 => x"2e098106",
   342 => x"86388053",
   343 => x"8ba304ff",
   344 => x"135372dd",
   345 => x"38868b2d",
   346 => x"9ce4089c",
   347 => x"f80c9ce4",
   348 => x"088b3881",
   349 => x"5287fc80",
   350 => x"d05183f1",
   351 => x"2d81ff0b",
   352 => x"d40c88bf",
   353 => x"2d9ce408",
   354 => x"9cfc0cd0",
   355 => x"08708f2a",
   356 => x"70810651",
   357 => x"515372f3",
   358 => x"3872d00c",
   359 => x"81ff0bd4",
   360 => x"0c815372",
   361 => x"9ce40c02",
   362 => x"8c050d04",
   363 => x"02f0050d",
   364 => x"805481ff",
   365 => x"0bd40cd0",
   366 => x"08708f2a",
   367 => x"70810651",
   368 => x"515372f3",
   369 => x"3882810b",
   370 => x"d00c81ff",
   371 => x"0bd40c75",
   372 => x"5287fc80",
   373 => x"d15183f1",
   374 => x"2d9ce408",
   375 => x"9e388480",
   376 => x"52765187",
   377 => x"b72d9ce4",
   378 => x"0854d008",
   379 => x"708f2a70",
   380 => x"81065151",
   381 => x"5372f338",
   382 => x"72d00c73",
   383 => x"9ce40c02",
   384 => x"90050d04",
   385 => x"02f4050d",
   386 => x"7470882a",
   387 => x"83fe8006",
   388 => x"7072982a",
   389 => x"0772882b",
   390 => x"87fc8080",
   391 => x"0673982b",
   392 => x"81f00a06",
   393 => x"71730707",
   394 => x"9ce40c56",
   395 => x"51535102",
   396 => x"8c050d04",
   397 => x"02f8050d",
   398 => x"028e0580",
   399 => x"f52d7488",
   400 => x"2b077083",
   401 => x"ffff069c",
   402 => x"e40c5102",
   403 => x"88050d04",
   404 => x"02f8050d",
   405 => x"7370902b",
   406 => x"71902a07",
   407 => x"9ce40c52",
   408 => x"0288050d",
   409 => x"0402f405",
   410 => x"0d9cf408",
   411 => x"53cc0870",
   412 => x"82800652",
   413 => x"5270732e",
   414 => x"f4387282",
   415 => x"80329cf4",
   416 => x"0c71fdff",
   417 => x"069ce40c",
   418 => x"028c050d",
   419 => x"0402f405",
   420 => x"0d800b9c",
   421 => x"f40c8ce5",
   422 => x"2d9ce408",
   423 => x"529cf408",
   424 => x"802e8638",
   425 => x"ad518dac",
   426 => x"0480df51",
   427 => x"81f72d71",
   428 => x"81812e80",
   429 => x"ec387181",
   430 => x"81248a38",
   431 => x"7181802e",
   432 => x"8d388ec9",
   433 => x"04718182",
   434 => x"2e93388e",
   435 => x"c90499f0",
   436 => x"5182bb2d",
   437 => x"9cf40872",
   438 => x"07528e9b",
   439 => x"0499fc51",
   440 => x"82bb2d9c",
   441 => x"fc0b80f5",
   442 => x"2d9cf408",
   443 => x"07cc0c8c",
   444 => x"e52d9cfd",
   445 => x"0b80f52d",
   446 => x"9cf40807",
   447 => x"cc0c8ce5",
   448 => x"2d9cfe0b",
   449 => x"80f52d9c",
   450 => x"f40807cc",
   451 => x"0c8ce52d",
   452 => x"9cff0b80",
   453 => x"f52d9cf4",
   454 => x"08075271",
   455 => x"cc0c8ecf",
   456 => x"049a9051",
   457 => x"82bb2dbf",
   458 => x"ff538383",
   459 => x"2d9ce408",
   460 => x"81ff0670",
   461 => x"9cf40807",
   462 => x"cc0c528c",
   463 => x"e52dff13",
   464 => x"53728025",
   465 => x"e5388ecf",
   466 => x"049aa051",
   467 => x"82bb2d9a",
   468 => x"b45182bb",
   469 => x"2d8d9604",
   470 => x"02fc050d",
   471 => x"9ad05182",
   472 => x"bb2d8a8a",
   473 => x"2d9ce408",
   474 => x"802ea338",
   475 => x"9ae85182",
   476 => x"bb2d8fd6",
   477 => x"2d9b8051",
   478 => x"8d8d2d9c",
   479 => x"e408802e",
   480 => x"87389b8c",
   481 => x"518f8b04",
   482 => x"9b985182",
   483 => x"bb2d800b",
   484 => x"9ce40c02",
   485 => x"84050d04",
   486 => x"02e8050d",
   487 => x"77797b58",
   488 => x"55558053",
   489 => x"727625a3",
   490 => x"38747081",
   491 => x"055680f5",
   492 => x"2d747081",
   493 => x"055680f5",
   494 => x"2d525271",
   495 => x"712e8638",
   496 => x"81518fcd",
   497 => x"04811353",
   498 => x"8fa40480",
   499 => x"51709ce4",
   500 => x"0c029805",
   501 => x"0d0402d8",
   502 => x"050d800b",
   503 => x"a1d00c9b",
   504 => x"ac5182bb",
   505 => x"2d9dac52",
   506 => x"80518bac",
   507 => x"2d9ce408",
   508 => x"549ce408",
   509 => x"8c389bbc",
   510 => x"5182bb2d",
   511 => x"73559583",
   512 => x"049bd051",
   513 => x"82bb2d80",
   514 => x"56810b9d",
   515 => x"a00c8853",
   516 => x"9be8529d",
   517 => x"e2518f98",
   518 => x"2d9ce408",
   519 => x"762e0981",
   520 => x"0687389c",
   521 => x"e4089da0",
   522 => x"0c88539b",
   523 => x"f4529dfe",
   524 => x"518f982d",
   525 => x"9ce40887",
   526 => x"389ce408",
   527 => x"9da00c9d",
   528 => x"a008802e",
   529 => x"80ff38a0",
   530 => x"f20b80f5",
   531 => x"2da0f30b",
   532 => x"80f52d71",
   533 => x"982b7190",
   534 => x"2b07a0f4",
   535 => x"0b80f52d",
   536 => x"70882b72",
   537 => x"07a0f50b",
   538 => x"80f52d71",
   539 => x"07a1aa0b",
   540 => x"80f52da1",
   541 => x"ab0b80f5",
   542 => x"2d71882b",
   543 => x"07535f54",
   544 => x"525a5657",
   545 => x"557381ab",
   546 => x"aa2e0981",
   547 => x"068d3875",
   548 => x"518c842d",
   549 => x"9ce40856",
   550 => x"91ab0473",
   551 => x"82d4d52e",
   552 => x"8a389c80",
   553 => x"5182bb2d",
   554 => x"92cf049d",
   555 => x"ac527551",
   556 => x"8bac2d9c",
   557 => x"e408559c",
   558 => x"e408802e",
   559 => x"83c5389c",
   560 => x"a05182bb",
   561 => x"2d88539b",
   562 => x"f4529dfe",
   563 => x"518f982d",
   564 => x"9ce40889",
   565 => x"38810ba1",
   566 => x"d00c91f5",
   567 => x"0488539b",
   568 => x"e8529de2",
   569 => x"518f982d",
   570 => x"80559ce4",
   571 => x"08752e09",
   572 => x"8106838f",
   573 => x"38a1aa0b",
   574 => x"80f52d54",
   575 => x"7380d52e",
   576 => x"09810680",
   577 => x"ca38a1ab",
   578 => x"0b80f52d",
   579 => x"547381aa",
   580 => x"2e098106",
   581 => x"ba38800b",
   582 => x"9dac0b80",
   583 => x"f52d5654",
   584 => x"7481e92e",
   585 => x"83388154",
   586 => x"7481eb2e",
   587 => x"8c388055",
   588 => x"73752e09",
   589 => x"810682cb",
   590 => x"389db70b",
   591 => x"80f52d55",
   592 => x"748d389d",
   593 => x"b80b80f5",
   594 => x"2d547382",
   595 => x"2e863880",
   596 => x"55958304",
   597 => x"9db90b80",
   598 => x"f52d70a1",
   599 => x"d80cff05",
   600 => x"a1cc0c9d",
   601 => x"ba0b80f5",
   602 => x"2d9dbb0b",
   603 => x"80f52d58",
   604 => x"76057782",
   605 => x"80290570",
   606 => x"a1c00c9d",
   607 => x"bc0b80f5",
   608 => x"2d70a1bc",
   609 => x"0ca1d008",
   610 => x"59575876",
   611 => x"802e81a3",
   612 => x"3888539b",
   613 => x"f4529dfe",
   614 => x"518f982d",
   615 => x"9ce40881",
   616 => x"e238a1d8",
   617 => x"0870842b",
   618 => x"a1ac0c70",
   619 => x"a1d40c9d",
   620 => x"d10b80f5",
   621 => x"2d9dd00b",
   622 => x"80f52d71",
   623 => x"82802905",
   624 => x"9dd20b80",
   625 => x"f52d7084",
   626 => x"80802912",
   627 => x"9dd30b80",
   628 => x"f52d7081",
   629 => x"800a2912",
   630 => x"709da40c",
   631 => x"a1bc0871",
   632 => x"29a1c008",
   633 => x"0570a1e0",
   634 => x"0c9dd90b",
   635 => x"80f52d9d",
   636 => x"d80b80f5",
   637 => x"2d718280",
   638 => x"29059dda",
   639 => x"0b80f52d",
   640 => x"70848080",
   641 => x"29129ddb",
   642 => x"0b80f52d",
   643 => x"70982b81",
   644 => x"f00a0672",
   645 => x"05709da8",
   646 => x"0cfe117e",
   647 => x"297705a1",
   648 => x"c80c5259",
   649 => x"5243545e",
   650 => x"51525952",
   651 => x"5d575957",
   652 => x"9581049d",
   653 => x"be0b80f5",
   654 => x"2d9dbd0b",
   655 => x"80f52d71",
   656 => x"82802905",
   657 => x"70a1ac0c",
   658 => x"70a02983",
   659 => x"ff057089",
   660 => x"2a70a1d4",
   661 => x"0c9dc30b",
   662 => x"80f52d9d",
   663 => x"c20b80f5",
   664 => x"2d718280",
   665 => x"2905709d",
   666 => x"a40c7b71",
   667 => x"291e70a1",
   668 => x"c80c7d9d",
   669 => x"a80c7305",
   670 => x"a1e00c55",
   671 => x"5e515155",
   672 => x"55815574",
   673 => x"9ce40c02",
   674 => x"a8050d04",
   675 => x"02ec050d",
   676 => x"7670872c",
   677 => x"7180ff06",
   678 => x"555654a1",
   679 => x"d0088a38",
   680 => x"73882c74",
   681 => x"81ff0654",
   682 => x"559dac52",
   683 => x"a1c00815",
   684 => x"518bac2d",
   685 => x"9ce40854",
   686 => x"9ce40880",
   687 => x"2eb338a1",
   688 => x"d008802e",
   689 => x"98387284",
   690 => x"299dac05",
   691 => x"70085253",
   692 => x"8c842d9c",
   693 => x"e408f00a",
   694 => x"065395ef",
   695 => x"0472109d",
   696 => x"ac057080",
   697 => x"e02d5253",
   698 => x"8cb42d9c",
   699 => x"e4085372",
   700 => x"54739ce4",
   701 => x"0c029405",
   702 => x"0d0402c8",
   703 => x"050d7f61",
   704 => x"5f5b800b",
   705 => x"9da808a1",
   706 => x"c808595d",
   707 => x"56a1d008",
   708 => x"762e8a38",
   709 => x"a1d80884",
   710 => x"2b5896a3",
   711 => x"04a1d408",
   712 => x"842b5880",
   713 => x"59787827",
   714 => x"81a93878",
   715 => x"8f06a017",
   716 => x"5754738f",
   717 => x"389dac52",
   718 => x"76518117",
   719 => x"578bac2d",
   720 => x"9dac5680",
   721 => x"7680f52d",
   722 => x"56547474",
   723 => x"2e833881",
   724 => x"547481e5",
   725 => x"2e80f638",
   726 => x"81707506",
   727 => x"555d7380",
   728 => x"2e80ea38",
   729 => x"8b1680f5",
   730 => x"2d98065a",
   731 => x"7980de38",
   732 => x"8b537d52",
   733 => x"75518f98",
   734 => x"2d9ce408",
   735 => x"80cf389c",
   736 => x"1608518c",
   737 => x"842d9ce4",
   738 => x"08841c0c",
   739 => x"9a1680e0",
   740 => x"2d518cb4",
   741 => x"2d9ce408",
   742 => x"9ce40888",
   743 => x"1d0c9ce4",
   744 => x"085555a1",
   745 => x"d008802e",
   746 => x"98389416",
   747 => x"80e02d51",
   748 => x"8cb42d9c",
   749 => x"e408902b",
   750 => x"83fff00a",
   751 => x"06701651",
   752 => x"5473881c",
   753 => x"0c797b0c",
   754 => x"7c549889",
   755 => x"04811959",
   756 => x"96a504a1",
   757 => x"d008802e",
   758 => x"ae387b51",
   759 => x"958c2d9c",
   760 => x"e4089ce4",
   761 => x"0880ffff",
   762 => x"fff80655",
   763 => x"5c7380ff",
   764 => x"fffff82e",
   765 => x"92389ce4",
   766 => x"08fe05a1",
   767 => x"d80829a1",
   768 => x"e0080557",
   769 => x"96a30480",
   770 => x"54739ce4",
   771 => x"0c02b805",
   772 => x"0d0402f4",
   773 => x"050d7470",
   774 => x"08810571",
   775 => x"0c7008a1",
   776 => x"cc080653",
   777 => x"53718e38",
   778 => x"88130851",
   779 => x"958c2d9c",
   780 => x"e4088814",
   781 => x"0c810b9c",
   782 => x"e40c028c",
   783 => x"050d0402",
   784 => x"f0050d75",
   785 => x"881108fe",
   786 => x"05a1d808",
   787 => x"29a1e008",
   788 => x"117208a1",
   789 => x"cc080605",
   790 => x"79555354",
   791 => x"548bac2d",
   792 => x"9ce40853",
   793 => x"9ce40880",
   794 => x"2e833881",
   795 => x"53729ce4",
   796 => x"0c029005",
   797 => x"0d0402ec",
   798 => x"050d7777",
   799 => x"53a1b052",
   800 => x"5395fa2d",
   801 => x"9ce40854",
   802 => x"9ce40880",
   803 => x"2ebf389c",
   804 => x"c85182bb",
   805 => x"2da1b408",
   806 => x"83ff0589",
   807 => x"2a558054",
   808 => x"737525a7",
   809 => x"387252a1",
   810 => x"b05198bf",
   811 => x"2d9ce408",
   812 => x"802e9138",
   813 => x"a1b05198",
   814 => x"922d8480",
   815 => x"13811555",
   816 => x"5399a004",
   817 => x"9ce40854",
   818 => x"99cd0481",
   819 => x"54739ce4",
   820 => x"0c029405",
   821 => x"0d040000",
   822 => x"00ffffff",
   823 => x"ff00ffff",
   824 => x"ffff00ff",
   825 => x"ffffff00",
   826 => x"434d4400",
   827 => x"53504900",
   828 => x"476f7420",
   829 => x"4e4f500a",
   830 => x"00000000",
   831 => x"476f7420",
   832 => x"52454144",
   833 => x"43415041",
   834 => x"43495459",
   835 => x"0a000000",
   836 => x"476f7420",
   837 => x"424f4f54",
   838 => x"53545241",
   839 => x"500a0000",
   840 => x"756e6b6e",
   841 => x"6f776e20",
   842 => x"636f6d6d",
   843 => x"616e640a",
   844 => x"00000000",
   845 => x"57616974",
   846 => x"696e6720",
   847 => x"666f7220",
   848 => x"6e657874",
   849 => x"20636f6d",
   850 => x"6d616e64",
   851 => x"0a000000",
   852 => x"496e6974",
   853 => x"69616c69",
   854 => x"7a696e67",
   855 => x"20534420",
   856 => x"63617264",
   857 => x"0a000000",
   858 => x"48756e74",
   859 => x"696e6720",
   860 => x"666f7220",
   861 => x"70617274",
   862 => x"6974696f",
   863 => x"6e0a0000",
   864 => x"42494f53",
   865 => x"4e455854",
   866 => x"31383600",
   867 => x"42494f53",
   868 => x"2053656e",
   869 => x"740a0000",
   870 => x"42494f53",
   871 => x"204c6f61",
   872 => x"64206661",
   873 => x"696c6564",
   874 => x"0a000000",
   875 => x"52656164",
   876 => x"696e6720",
   877 => x"4d42520a",
   878 => x"00000000",
   879 => x"52656164",
   880 => x"206f6620",
   881 => x"4d425220",
   882 => x"6661696c",
   883 => x"65640a00",
   884 => x"4d425220",
   885 => x"73756363",
   886 => x"65737366",
   887 => x"756c6c79",
   888 => x"20726561",
   889 => x"640a0000",
   890 => x"46415431",
   891 => x"36202020",
   892 => x"00000000",
   893 => x"46415433",
   894 => x"32202020",
   895 => x"00000000",
   896 => x"4e6f2070",
   897 => x"61727469",
   898 => x"74696f6e",
   899 => x"20736967",
   900 => x"6e617475",
   901 => x"72652066",
   902 => x"6f756e64",
   903 => x"0a000000",
   904 => x"52656164",
   905 => x"20626f6f",
   906 => x"74207365",
   907 => x"63746f72",
   908 => x"2066726f",
   909 => x"6d206669",
   910 => x"72737420",
   911 => x"70617274",
   912 => x"6974696f",
   913 => x"6e0a0000",
   914 => x"4f70656e",
   915 => x"65642066",
   916 => x"696c652c",
   917 => x"206c6f61",
   918 => x"64696e67",
   919 => x"2e2e2e0a",
   920 => x"002e2e0a",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;


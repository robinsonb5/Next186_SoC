-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Bootstrap_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Bootstrap_ROM1;

architecture arch of Bootstrap_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0ba5",
     9 => x"d0080b0b",
    10 => x"0ba5d408",
    11 => x"0b0b0ba5",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a5d80c0b",
    16 => x"0b0ba5d4",
    17 => x"0c0b0b0b",
    18 => x"a5d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba38c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a5d070ab",
    57 => x"a4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8fd00402",
    62 => x"ec050d76",
    63 => x"53805572",
    64 => x"752e80c7",
    65 => x"38875472",
    66 => x"9c2a7384",
    67 => x"2b545271",
    68 => x"802e8338",
    69 => x"81558972",
    70 => x"259938b7",
    71 => x"1252749b",
    72 => x"38ff1454",
    73 => x"738025df",
    74 => x"38800ba5",
    75 => x"d00c0294",
    76 => x"050d04b0",
    77 => x"12527480",
    78 => x"2ee73871",
    79 => x"5182da2d",
    80 => x"ff145473",
    81 => x"8025c038",
    82 => x"82a904b0",
    83 => x"5182da2d",
    84 => x"800ba5d0",
    85 => x"0c029405",
    86 => x"0d0402f8",
    87 => x"050d7352",
    88 => x"c0087088",
    89 => x"2a708106",
    90 => x"51515170",
    91 => x"802ef138",
    92 => x"71c00c71",
    93 => x"a5d00c02",
    94 => x"88050d04",
    95 => x"02f8050d",
    96 => x"7352c408",
    97 => x"70882a70",
    98 => x"81065151",
    99 => x"5170802e",
   100 => x"f13871c4",
   101 => x"0c71a5d0",
   102 => x"0c028805",
   103 => x"0d0402e8",
   104 => x"050d8078",
   105 => x"57557570",
   106 => x"84055708",
   107 => x"53805472",
   108 => x"982a7388",
   109 => x"2b545271",
   110 => x"802ea238",
   111 => x"c0087088",
   112 => x"2a708106",
   113 => x"51515170",
   114 => x"802ef138",
   115 => x"71c00c81",
   116 => x"15811555",
   117 => x"55837425",
   118 => x"d63871ca",
   119 => x"3874a5d0",
   120 => x"0c029805",
   121 => x"0d0402f4",
   122 => x"050dd452",
   123 => x"81ff720c",
   124 => x"71085381",
   125 => x"ff720c72",
   126 => x"882b83fe",
   127 => x"80067208",
   128 => x"7081ff06",
   129 => x"51525381",
   130 => x"ff720c72",
   131 => x"7107882b",
   132 => x"72087081",
   133 => x"ff065152",
   134 => x"5381ff72",
   135 => x"0c727107",
   136 => x"882b7208",
   137 => x"7081ff06",
   138 => x"7207a5d0",
   139 => x"0c525302",
   140 => x"8c050d04",
   141 => x"02f4050d",
   142 => x"74767181",
   143 => x"ff06d40c",
   144 => x"5353a6b4",
   145 => x"08853871",
   146 => x"892b5271",
   147 => x"982ad40c",
   148 => x"71902a70",
   149 => x"81ff06d4",
   150 => x"0c517188",
   151 => x"2a7081ff",
   152 => x"06d40c51",
   153 => x"7181ff06",
   154 => x"d40c7290",
   155 => x"2a7081ff",
   156 => x"06d40c51",
   157 => x"d4087081",
   158 => x"ff065151",
   159 => x"82b8bf52",
   160 => x"7081ff2e",
   161 => x"09810694",
   162 => x"3881ff0b",
   163 => x"d40cd408",
   164 => x"7081ff06",
   165 => x"ff145451",
   166 => x"5171e538",
   167 => x"70a5d00c",
   168 => x"028c050d",
   169 => x"0402fc05",
   170 => x"0d81c751",
   171 => x"81ff0bd4",
   172 => x"0cff1151",
   173 => x"708025f4",
   174 => x"38028405",
   175 => x"0d0402f0",
   176 => x"050d85a5",
   177 => x"2d819c9f",
   178 => x"53805287",
   179 => x"fc80f751",
   180 => x"84b42da5",
   181 => x"d00854a5",
   182 => x"d008812e",
   183 => x"9038ff13",
   184 => x"5372e638",
   185 => x"72a5d00c",
   186 => x"0290050d",
   187 => x"0481ff0b",
   188 => x"d40c820a",
   189 => x"52849c80",
   190 => x"e95184b4",
   191 => x"2da5d008",
   192 => x"802e8e38",
   193 => x"85a52dff",
   194 => x"135372ff",
   195 => x"bc3885e4",
   196 => x"0481ff0b",
   197 => x"d40c73a5",
   198 => x"d00c0290",
   199 => x"050d0402",
   200 => x"f4050d81",
   201 => x"ff0bd40c",
   202 => x"a39c5183",
   203 => x"9e2d9353",
   204 => x"805287fc",
   205 => x"80c15184",
   206 => x"b42da5d0",
   207 => x"08802e93",
   208 => x"3885a52d",
   209 => x"ff135372",
   210 => x"e73872a5",
   211 => x"d00c028c",
   212 => x"050d0481",
   213 => x"ff0bd40c",
   214 => x"810ba5d0",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050d85a5",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"5184b42d",
   221 => x"a5d00881",
   222 => x"2e8f3886",
   223 => x"9f2d8054",
   224 => x"73a5d00c",
   225 => x"0290050d",
   226 => x"0483e62d",
   227 => x"a5d00883",
   228 => x"ffff0653",
   229 => x"7283aa2e",
   230 => x"098106df",
   231 => x"3881ff0b",
   232 => x"d40cb153",
   233 => x"85be2da5",
   234 => x"d0089538",
   235 => x"72822ece",
   236 => x"38ff1353",
   237 => x"72ee3872",
   238 => x"a5d00c02",
   239 => x"90050d04",
   240 => x"805287fc",
   241 => x"80fa5184",
   242 => x"b42da5d0",
   243 => x"08de3881",
   244 => x"ff0bd40c",
   245 => x"d4085381",
   246 => x"ff0bd40c",
   247 => x"81ff0bd4",
   248 => x"0c81ff0b",
   249 => x"d40c81ff",
   250 => x"0bd40c72",
   251 => x"862a7081",
   252 => x"06a5d008",
   253 => x"56515372",
   254 => x"802eff84",
   255 => x"38810ba5",
   256 => x"d00c0290",
   257 => x"050d0402",
   258 => x"e8050d78",
   259 => x"5681ff0b",
   260 => x"d40cd008",
   261 => x"708f2a70",
   262 => x"81065151",
   263 => x"5372f338",
   264 => x"82810bd0",
   265 => x"0c81ff0b",
   266 => x"d40c7752",
   267 => x"87fc80d8",
   268 => x"5184b42d",
   269 => x"a5d00881",
   270 => x"823881ff",
   271 => x"0bd40c81",
   272 => x"fe0bd40c",
   273 => x"80ff5575",
   274 => x"70840557",
   275 => x"0870982a",
   276 => x"d40c7090",
   277 => x"2c7081ff",
   278 => x"06d40c54",
   279 => x"70882c70",
   280 => x"81ff06d4",
   281 => x"0c547081",
   282 => x"ff06d40c",
   283 => x"54ff1555",
   284 => x"748025d3",
   285 => x"3881ff0b",
   286 => x"d40c81ff",
   287 => x"0bd40c81",
   288 => x"ff0bd40c",
   289 => x"868da054",
   290 => x"81ff0bd4",
   291 => x"0cd40881",
   292 => x"ff065574",
   293 => x"8738ff14",
   294 => x"5473ed38",
   295 => x"81ff0bd4",
   296 => x"0cd00870",
   297 => x"8f2a7081",
   298 => x"06515153",
   299 => x"72f33872",
   300 => x"d00c72a5",
   301 => x"d00c0298",
   302 => x"050d04a3",
   303 => x"a051839e",
   304 => x"2d810ba5",
   305 => x"d00c0298",
   306 => x"050d0402",
   307 => x"ec050d76",
   308 => x"78545480",
   309 => x"5580dbc6",
   310 => x"df5281ff",
   311 => x"0bd40cd4",
   312 => x"087081ff",
   313 => x"06515170",
   314 => x"81fe2e95",
   315 => x"38ff1252",
   316 => x"71e83881",
   317 => x"ff0bd40c",
   318 => x"74a5d00c",
   319 => x"0294050d",
   320 => x"04800ba6",
   321 => x"d80c8373",
   322 => x"259f3883",
   323 => x"e62da5d0",
   324 => x"08747084",
   325 => x"05560ca6",
   326 => x"d808a5d0",
   327 => x"0805a6d8",
   328 => x"0cfc1353",
   329 => x"728324e3",
   330 => x"38807325",
   331 => x"a03881ff",
   332 => x"0bd40cff",
   333 => x"74708105",
   334 => x"5681b72d",
   335 => x"a6d80881",
   336 => x"ff05a6d8",
   337 => x"0cff1353",
   338 => x"728024e2",
   339 => x"38815581",
   340 => x"ff0bd40c",
   341 => x"74a5d00c",
   342 => x"0294050d",
   343 => x"0402e805",
   344 => x"0d805287",
   345 => x"fc80c951",
   346 => x"84b42d92",
   347 => x"52a6c451",
   348 => x"89cb2da6",
   349 => x"c40b80f5",
   350 => x"2d81c006",
   351 => x"537280c0",
   352 => x"2e80f738",
   353 => x"a6cd0b80",
   354 => x"f52d7010",
   355 => x"8606a6ce",
   356 => x"0b80f52d",
   357 => x"70872a72",
   358 => x"07a6c90b",
   359 => x"80f52d8f",
   360 => x"06a6ca0b",
   361 => x"80f52d70",
   362 => x"8a2b9880",
   363 => x"06a6cb0b",
   364 => x"80f52d70",
   365 => x"822b7207",
   366 => x"a6cc0b80",
   367 => x"f52d7086",
   368 => x"2a720782",
   369 => x"1881782b",
   370 => x"81138173",
   371 => x"2b712951",
   372 => x"53585852",
   373 => x"52525259",
   374 => x"53545258",
   375 => x"55558480",
   376 => x"75258e38",
   377 => x"72107581",
   378 => x"2c565374",
   379 => x"848024f4",
   380 => x"3872a5d0",
   381 => x"0c029805",
   382 => x"0d04a6cb",
   383 => x"0b80f52d",
   384 => x"a6cc0b80",
   385 => x"f52d7190",
   386 => x"2b71882b",
   387 => x"07a6cd0b",
   388 => x"80f52d71",
   389 => x"81fffe80",
   390 => x"06077088",
   391 => x"80298880",
   392 => x"05a5d00c",
   393 => x"51555755",
   394 => x"0298050d",
   395 => x"0402f405",
   396 => x"0d810ba6",
   397 => x"b40cd008",
   398 => x"708f2a70",
   399 => x"81065151",
   400 => x"5372f338",
   401 => x"72d00c85",
   402 => x"a52da3b0",
   403 => x"51839e2d",
   404 => x"d008708f",
   405 => x"2a708106",
   406 => x"51515372",
   407 => x"f338810b",
   408 => x"d00c8753",
   409 => x"805284d4",
   410 => x"80c05184",
   411 => x"b42da5d0",
   412 => x"08812e8d",
   413 => x"3872822e",
   414 => x"80c538ff",
   415 => x"135372e4",
   416 => x"3886e22d",
   417 => x"a5d008a6",
   418 => x"b40ca5d0",
   419 => x"08802eb9",
   420 => x"3881ff0b",
   421 => x"d40c8add",
   422 => x"2da5d008",
   423 => x"a6b80cd0",
   424 => x"08708f2a",
   425 => x"70810651",
   426 => x"515372f3",
   427 => x"3872d00c",
   428 => x"81ff0bd4",
   429 => x"0c810ba5",
   430 => x"d00c028c",
   431 => x"050d0480",
   432 => x"0ba5d00c",
   433 => x"028c050d",
   434 => x"04815287",
   435 => x"fc80d051",
   436 => x"84b42d81",
   437 => x"ff0bd40c",
   438 => x"8add2da5",
   439 => x"d008a6b8",
   440 => x"0c8d9f04",
   441 => x"02f0050d",
   442 => x"805481ff",
   443 => x"0bd40cd0",
   444 => x"08708f2a",
   445 => x"70810651",
   446 => x"515372f3",
   447 => x"3882810b",
   448 => x"d00c81ff",
   449 => x"0bd40c75",
   450 => x"5287fc80",
   451 => x"d15184b4",
   452 => x"2da5d008",
   453 => x"802e8a38",
   454 => x"73a5d00c",
   455 => x"0290050d",
   456 => x"04848052",
   457 => x"765189cb",
   458 => x"2da5d008",
   459 => x"54d00870",
   460 => x"8f2a7081",
   461 => x"06515153",
   462 => x"72f33872",
   463 => x"d00c73a5",
   464 => x"d00c0290",
   465 => x"050d0402",
   466 => x"f4050d74",
   467 => x"70882a83",
   468 => x"fe800670",
   469 => x"72982a07",
   470 => x"72882b87",
   471 => x"fc808006",
   472 => x"73982b81",
   473 => x"f00a0671",
   474 => x"730707a5",
   475 => x"d00c5651",
   476 => x"5351028c",
   477 => x"050d0402",
   478 => x"f8050d02",
   479 => x"8e0580f5",
   480 => x"2d74882b",
   481 => x"077083ff",
   482 => x"ff06a5d0",
   483 => x"0c510288",
   484 => x"050d0402",
   485 => x"f8050d73",
   486 => x"70902b71",
   487 => x"902a07a5",
   488 => x"d00c5202",
   489 => x"88050d04",
   490 => x"02f4050d",
   491 => x"a6b00853",
   492 => x"cc087082",
   493 => x"80065252",
   494 => x"70732ef4",
   495 => x"38728280",
   496 => x"32a6b00c",
   497 => x"71fdff06",
   498 => x"a5d00c02",
   499 => x"8c050d04",
   500 => x"02d8050d",
   501 => x"800ba6b0",
   502 => x"0ca3b451",
   503 => x"839e2d8c",
   504 => x"ad2d8054",
   505 => x"a5d00874",
   506 => x"2e098106",
   507 => x"8a3873a5",
   508 => x"d00c02a8",
   509 => x"050d04a3",
   510 => x"bc51839e",
   511 => x"2d97e92d",
   512 => x"8fa82da5",
   513 => x"d0085aa5",
   514 => x"d0088183",
   515 => x"2ebd38a5",
   516 => x"d0088183",
   517 => x"2482d838",
   518 => x"a5d00881",
   519 => x"812e838b",
   520 => x"38a5d008",
   521 => x"81812484",
   522 => x"a738a5d0",
   523 => x"0881802e",
   524 => x"86b438a3",
   525 => x"c451839e",
   526 => x"2d8fa82d",
   527 => x"a5d0085a",
   528 => x"a5d00881",
   529 => x"832e0981",
   530 => x"06c538a6",
   531 => x"b008cc0c",
   532 => x"8fa82da5",
   533 => x"d008982b",
   534 => x"a6b008cc",
   535 => x"0c588fa8",
   536 => x"2da5d008",
   537 => x"902b7807",
   538 => x"a6b008cc",
   539 => x"0c588fa8",
   540 => x"2da5d008",
   541 => x"882b7807",
   542 => x"a6b008cc",
   543 => x"0c588fa8",
   544 => x"2d77a5d0",
   545 => x"0807a6b0",
   546 => x"08cc0c58",
   547 => x"8fa82da5",
   548 => x"d0085990",
   549 => x"53805277",
   550 => x"5181f72d",
   551 => x"ff195978",
   552 => x"ff2e81c3",
   553 => x"38a6e857",
   554 => x"7981852e",
   555 => x"85c938a3",
   556 => x"cc51839e",
   557 => x"2d765277",
   558 => x"51811858",
   559 => x"8de42d80",
   560 => x"ff567670",
   561 => x"84055808",
   562 => x"70982aa6",
   563 => x"b00807cc",
   564 => x"0c558fa8",
   565 => x"2d74902a",
   566 => x"7081ff06",
   567 => x"70a6b008",
   568 => x"07cc0c51",
   569 => x"548fa82d",
   570 => x"74882a70",
   571 => x"81ff0670",
   572 => x"a6b00807",
   573 => x"cc0c5154",
   574 => x"8fa82d74",
   575 => x"81ff0670",
   576 => x"a6b00807",
   577 => x"cc0c558f",
   578 => x"a82dff16",
   579 => x"56807624",
   580 => x"ff8a3876",
   581 => x"70840558",
   582 => x"0870982a",
   583 => x"a6b00807",
   584 => x"cc0c558f",
   585 => x"a82d7490",
   586 => x"2a7081ff",
   587 => x"0670a6b0",
   588 => x"0807cc0c",
   589 => x"51548fa8",
   590 => x"2d74882a",
   591 => x"7081ff06",
   592 => x"70a6b008",
   593 => x"07cc0c51",
   594 => x"548fa82d",
   595 => x"7481ff06",
   596 => x"70a6b008",
   597 => x"07cc0c55",
   598 => x"8fa82dff",
   599 => x"16567580",
   600 => x"25fedf38",
   601 => x"919c04a6",
   602 => x"b008cc0c",
   603 => x"908004a5",
   604 => x"d0088185",
   605 => x"2efdd438",
   606 => x"81850ba5",
   607 => x"d0082482",
   608 => x"9a38a5d0",
   609 => x"0881fe2e",
   610 => x"098106fd",
   611 => x"a638a6b0",
   612 => x"0881fe07",
   613 => x"cc0c8fa8",
   614 => x"2da5d008",
   615 => x"5182da2d",
   616 => x"a6b00881",
   617 => x"fe07cc0c",
   618 => x"908004a3",
   619 => x"d051839e",
   620 => x"2da3d852",
   621 => x"aaec519e",
   622 => x"982da5d0",
   623 => x"0854a5d0",
   624 => x"08802e83",
   625 => x"ce38aaf0",
   626 => x"0883ff05",
   627 => x"892a5780",
   628 => x"55747725",
   629 => x"fcaa38a6",
   630 => x"e852aaec",
   631 => x"51a18f2d",
   632 => x"a5d00880",
   633 => x"2e80cb38",
   634 => x"a3e45183",
   635 => x"9e2d8056",
   636 => x"a6e81680",
   637 => x"f52da6b0",
   638 => x"0807cc0c",
   639 => x"8fa82da6",
   640 => x"b008802e",
   641 => x"b838ad51",
   642 => x"82da2d81",
   643 => x"165683ff",
   644 => x"7625dd38",
   645 => x"81155574",
   646 => x"7725fbe4",
   647 => x"38aaec51",
   648 => x"a0d62da6",
   649 => x"e852aaec",
   650 => x"51a18f2d",
   651 => x"a5d008ff",
   652 => x"b738a5d0",
   653 => x"08a5d00c",
   654 => x"02a8050d",
   655 => x"0480df51",
   656 => x"82da2d81",
   657 => x"165683ff",
   658 => x"7625ffa4",
   659 => x"38949404",
   660 => x"a3e85183",
   661 => x"9e2da3f0",
   662 => x"52aaec51",
   663 => x"9e982da6",
   664 => x"b80b80f5",
   665 => x"2da6b008",
   666 => x"07cc0c8f",
   667 => x"a82da6b9",
   668 => x"0b80f52d",
   669 => x"a6b00807",
   670 => x"cc0c8fa8",
   671 => x"2da6ba0b",
   672 => x"80f52da6",
   673 => x"b00807cc",
   674 => x"0c8fa82d",
   675 => x"a6bb0b80",
   676 => x"f52da6b0",
   677 => x"0807cc0c",
   678 => x"908004a3",
   679 => x"fc51839e",
   680 => x"2da6b008",
   681 => x"cc0c8fa8",
   682 => x"2da5d008",
   683 => x"982ba6b0",
   684 => x"08cc0c58",
   685 => x"8fa82da5",
   686 => x"d008902b",
   687 => x"7807a6b0",
   688 => x"08cc0c58",
   689 => x"8fa82da5",
   690 => x"d008882b",
   691 => x"7807a6b0",
   692 => x"08cc0c58",
   693 => x"8fa82d77",
   694 => x"a5d00807",
   695 => x"a6b008cc",
   696 => x"0c588fa8",
   697 => x"2da5d008",
   698 => x"59905380",
   699 => x"52775181",
   700 => x"f72dff19",
   701 => x"5978ff2e",
   702 => x"fced38a6",
   703 => x"e80ba480",
   704 => x"5255839e",
   705 => x"2d80ff56",
   706 => x"a6b008cc",
   707 => x"0c8fa82d",
   708 => x"a6b008cc",
   709 => x"0ca5d008",
   710 => x"882b548f",
   711 => x"a82da6b0",
   712 => x"08cc0c73",
   713 => x"a5d00807",
   714 => x"882b548f",
   715 => x"a82da6b0",
   716 => x"08cc0c73",
   717 => x"a5d00807",
   718 => x"882b548f",
   719 => x"a82d73a5",
   720 => x"d0080775",
   721 => x"70840557",
   722 => x"0cff1656",
   723 => x"758025ff",
   724 => x"b738a480",
   725 => x"51839e2d",
   726 => x"a6e85277",
   727 => x"51811858",
   728 => x"88872d95",
   729 => x"f204a484",
   730 => x"51839e2d",
   731 => x"a6b00881",
   732 => x"8007cc0c",
   733 => x"908004a4",
   734 => x"8c51839e",
   735 => x"2d7752aa",
   736 => x"ec51a1c6",
   737 => x"2d7652aa",
   738 => x"ec51a18f",
   739 => x"2d80ff56",
   740 => x"91c204a4",
   741 => x"9051839e",
   742 => x"2d73a5d0",
   743 => x"0c02a805",
   744 => x"0d0402e8",
   745 => x"050d7779",
   746 => x"7b585555",
   747 => x"80537276",
   748 => x"25a33874",
   749 => x"70810556",
   750 => x"80f52d74",
   751 => x"70810556",
   752 => x"80f52d52",
   753 => x"5271712e",
   754 => x"09810693",
   755 => x"38811353",
   756 => x"757324df",
   757 => x"38800ba5",
   758 => x"d00c0298",
   759 => x"050d0481",
   760 => x"0ba5d00c",
   761 => x"0298050d",
   762 => x"0402d805",
   763 => x"0d800bab",
   764 => x"900ca498",
   765 => x"51839e2d",
   766 => x"a6e85280",
   767 => x"518de42d",
   768 => x"a5d00854",
   769 => x"a5d00892",
   770 => x"38a4a851",
   771 => x"839e2d73",
   772 => x"5675a5d0",
   773 => x"0c02a805",
   774 => x"0d04a4bc",
   775 => x"51839e2d",
   776 => x"8055810b",
   777 => x"a6dc0c88",
   778 => x"53a4d452",
   779 => x"a79e5197",
   780 => x"a22da5d0",
   781 => x"08752e80",
   782 => x"fb388853",
   783 => x"a4e052a7",
   784 => x"ba5197a2",
   785 => x"2da5d008",
   786 => x"8738a5d0",
   787 => x"08a6dc0c",
   788 => x"a6dc0880",
   789 => x"2e818938",
   790 => x"aaae0b80",
   791 => x"f52daaaf",
   792 => x"0b80f52d",
   793 => x"71982b71",
   794 => x"902b07aa",
   795 => x"b00b80f5",
   796 => x"2d70882b",
   797 => x"7207aab1",
   798 => x"0b80f52d",
   799 => x"7107aae6",
   800 => x"0b80f52d",
   801 => x"aae70b80",
   802 => x"f52d7188",
   803 => x"2b075340",
   804 => x"55525a56",
   805 => x"57557381",
   806 => x"abaa2ea1",
   807 => x"387382d4",
   808 => x"d52ea338",
   809 => x"a4ec5183",
   810 => x"9e2d800b",
   811 => x"a5d00c02",
   812 => x"a8050d04",
   813 => x"a5d008a6",
   814 => x"dc0c98ba",
   815 => x"0474518e",
   816 => x"c72da5d0",
   817 => x"0855a6e8",
   818 => x"5274518d",
   819 => x"e42da5d0",
   820 => x"0856a5d0",
   821 => x"08802efe",
   822 => x"b838a58c",
   823 => x"51839e2d",
   824 => x"8853a4e0",
   825 => x"52a7ba51",
   826 => x"97a22da5",
   827 => x"d00881fa",
   828 => x"38810bab",
   829 => x"900caae6",
   830 => x"0b80f52d",
   831 => x"547380d5",
   832 => x"2e098106",
   833 => x"ffa438aa",
   834 => x"e70b80f5",
   835 => x"2d547381",
   836 => x"aa2e0981",
   837 => x"06ff9338",
   838 => x"800ba6e8",
   839 => x"0b80f52d",
   840 => x"57547581",
   841 => x"e92e8338",
   842 => x"81547581",
   843 => x"eb2e8c38",
   844 => x"80567376",
   845 => x"2e098106",
   846 => x"fdd738a6",
   847 => x"f30b80f5",
   848 => x"2d5675fe",
   849 => x"e538a6f4",
   850 => x"0b80f52d",
   851 => x"5473822e",
   852 => x"098106fe",
   853 => x"d538a6f5",
   854 => x"0b80f52d",
   855 => x"70ab980c",
   856 => x"ff05ab8c",
   857 => x"0ca6f60b",
   858 => x"80f52da6",
   859 => x"f70b80f5",
   860 => x"2d5b7505",
   861 => x"7a828029",
   862 => x"0570ab80",
   863 => x"0ca6f80b",
   864 => x"80f52d70",
   865 => x"aafc0cab",
   866 => x"90085b59",
   867 => x"577880f8",
   868 => x"38a6fa0b",
   869 => x"80f52da6",
   870 => x"f90b80f5",
   871 => x"2d718280",
   872 => x"290570aa",
   873 => x"e80c70a0",
   874 => x"2983ff05",
   875 => x"70892a70",
   876 => x"ab940ca6",
   877 => x"ff0b80f5",
   878 => x"2da6fe0b",
   879 => x"80f52d71",
   880 => x"82802905",
   881 => x"70a6e00c",
   882 => x"7d71291d",
   883 => x"70ab880c",
   884 => x"7fa6e40c",
   885 => x"7305aba0",
   886 => x"0c5a5a51",
   887 => x"51555a81",
   888 => x"5675a5d0",
   889 => x"0c02a805",
   890 => x"0d048853",
   891 => x"a4d452a7",
   892 => x"9e5197a2",
   893 => x"2d8056a5",
   894 => x"d008762e",
   895 => x"fdf83875",
   896 => x"a5d00c02",
   897 => x"a8050d04",
   898 => x"8853a4e0",
   899 => x"52a7ba51",
   900 => x"97a22da5",
   901 => x"d008fbf9",
   902 => x"38ab9808",
   903 => x"70842baa",
   904 => x"e80c70ab",
   905 => x"940ca78d",
   906 => x"0b80f52d",
   907 => x"a78c0b80",
   908 => x"f52d7182",
   909 => x"802905a7",
   910 => x"8e0b80f5",
   911 => x"2d708480",
   912 => x"802912a7",
   913 => x"8f0b80f5",
   914 => x"2d708180",
   915 => x"0a291270",
   916 => x"a6e00caa",
   917 => x"fc087129",
   918 => x"ab800805",
   919 => x"70aba00c",
   920 => x"a7950b80",
   921 => x"f52da794",
   922 => x"0b80f52d",
   923 => x"71828029",
   924 => x"05a7960b",
   925 => x"80f52d70",
   926 => x"84808029",
   927 => x"12a7970b",
   928 => x"80f52d70",
   929 => x"982b81f0",
   930 => x"0a067205",
   931 => x"70a6e40c",
   932 => x"fe117e29",
   933 => x"7705ab88",
   934 => x"0c525952",
   935 => x"55585e51",
   936 => x"525f525b",
   937 => x"57555781",
   938 => x"569be104",
   939 => x"02ec050d",
   940 => x"7670872c",
   941 => x"7180ff06",
   942 => x"565653ab",
   943 => x"90088a38",
   944 => x"72882c73",
   945 => x"81ff0655",
   946 => x"55a6e852",
   947 => x"ab800815",
   948 => x"518de42d",
   949 => x"a5d00853",
   950 => x"a5d00880",
   951 => x"2e9c38ab",
   952 => x"9008802e",
   953 => x"9e387310",
   954 => x"10a6e805",
   955 => x"70085253",
   956 => x"8ec72da5",
   957 => x"d008f00a",
   958 => x"065372a5",
   959 => x"d00c0294",
   960 => x"050d0473",
   961 => x"10a6e805",
   962 => x"7080e02d",
   963 => x"52538ef7",
   964 => x"2da5d008",
   965 => x"539dfa04",
   966 => x"02cc050d",
   967 => x"7e605d5d",
   968 => x"800ba6e4",
   969 => x"08ab8808",
   970 => x"5a5c57ab",
   971 => x"9008772e",
   972 => x"818a38ab",
   973 => x"9808842b",
   974 => x"59805675",
   975 => x"792780c4",
   976 => x"38758f06",
   977 => x"a0185854",
   978 => x"73802e80",
   979 => x"fa388077",
   980 => x"80f52d55",
   981 => x"5573752e",
   982 => x"83388155",
   983 => x"7381e52e",
   984 => x"9a388170",
   985 => x"7606555a",
   986 => x"73802e8f",
   987 => x"388b1780",
   988 => x"f52d9806",
   989 => x"5574802e",
   990 => x"80de3881",
   991 => x"16567876",
   992 => x"26ffbe38",
   993 => x"ab900880",
   994 => x"2e81c138",
   995 => x"7a519dac",
   996 => x"2da5d008",
   997 => x"a5d00880",
   998 => x"fffffff8",
   999 => x"06555b73",
  1000 => x"80ffffff",
  1001 => x"f82e81a4",
  1002 => x"38a5d008",
  1003 => x"fe05ab98",
  1004 => x"0829aba0",
  1005 => x"08055880",
  1006 => x"569ebb04",
  1007 => x"ab940884",
  1008 => x"2b598056",
  1009 => x"9ebb04a6",
  1010 => x"e8527751",
  1011 => x"8118588d",
  1012 => x"e42da6e8",
  1013 => x"579ece04",
  1014 => x"8b537b52",
  1015 => x"765197a2",
  1016 => x"2da5d008",
  1017 => x"ff95389c",
  1018 => x"1708518e",
  1019 => x"c72da5d0",
  1020 => x"08841e0c",
  1021 => x"9a1780e0",
  1022 => x"2d518ef7",
  1023 => x"2da5d008",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

